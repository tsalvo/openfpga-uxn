-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity inc2_0CLK_263c9bc8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_263c9bc8;
architecture arch of inc2_0CLK_263c9bc8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1327_c6_2b9e]
signal BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1327_c2_a117]
signal t16_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1327_c2_a117]
signal tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1327_c2_a117]
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1327_c2_a117]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1327_c2_a117]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1327_c2_a117]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1327_c2_a117]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1334_c11_f617]
signal BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal t16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1334_c7_e39f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1337_c11_1951]
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal t16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1337_c7_15c1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l1339_c3_8499]
signal CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1341_c11_a89f]
signal BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1341_c7_d4b7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1342_c3_f5e1]
signal BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1343_c11_3ebf]
signal BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output : unsigned(16 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1345_c30_bd88]
signal sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1350_c11_03f4]
signal BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1350_c7_6af6]
signal result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1350_c7_6af6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1350_c7_6af6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1350_c7_6af6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1350_c7_6af6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : signed(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l1353_c31_f4c2]
signal CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1355_c11_e864]
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c7_a636]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c7_a636]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e
BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_left,
BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_right,
BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output);

-- t16_MUX_uxn_opcodes_h_l1327_c2_a117
t16_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
t16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
t16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1327_c2_a117
tmp16_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117
result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_left,
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_right,
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output);

-- t16_MUX_uxn_opcodes_h_l1334_c7_e39f
t16_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f
tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_left,
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_right,
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output);

-- t16_MUX_uxn_opcodes_h_l1337_c7_15c1
t16_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1
tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1
result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output);

-- CONST_SL_8_uxn_opcodes_h_l1339_c3_8499
CONST_SL_8_uxn_opcodes_h_l1339_c3_8499 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_x,
CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_left,
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_right,
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output);

-- t16_MUX_uxn_opcodes_h_l1341_c7_d4b7
t16_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7
tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7
result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1
BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_left,
BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_right,
BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf
BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_left,
BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_right,
BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88
sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_ins,
sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_x,
sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_y,
sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4
BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_left,
BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_right,
BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6
result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6
result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6
result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output);

-- CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2
CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_x,
CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864
BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_left,
BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_right,
BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output,
 t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output,
 t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output,
 t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output,
 CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output,
 t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output,
 sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output,
 CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1331_c3_a5a8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1335_c3_1c1d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_uxn_opcodes_h_l1343_c3_1378 : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1347_c3_030f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output : unsigned(16 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1348_c21_f3c2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1352_c3_722e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1351_c3_2327 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1353_c21_ff03_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1338_l1342_DUPLICATE_cb7b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1350_l1337_DUPLICATE_8ec4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1323_l1360_DUPLICATE_ca38_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1352_c3_722e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1352_c3_722e;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1347_c3_030f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1347_c3_030f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1331_c3_a5a8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1331_c3_a5a8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1335_c3_1c1d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1335_c3_1c1d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1351_c3_2327 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1351_c3_2327;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := tmp16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1345_c30_bd88] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_ins;
     sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_x;
     sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output := sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1350_l1337_DUPLICATE_8ec4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1350_l1337_DUPLICATE_8ec4_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1334_c11_f617] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_left;
     BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output := BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1350_c11_03f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1338_l1342_DUPLICATE_cb7b LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1338_l1342_DUPLICATE_cb7b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1341_c11_a89f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l1353_c31_f4c2] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_x <= VAR_CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output := CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1327_c6_2b9e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1355_c11_e864] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_left;
     BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output := BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1337_c11_1951] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_left;
     BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output := BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c6_2b9e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_f617_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_1951_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_a89f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1350_c11_03f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c11_e864_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1338_l1342_DUPLICATE_cb7b_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1338_l1342_DUPLICATE_cb7b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_f715_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1350_l1341_l1337_l1355_l1334_DUPLICATE_4b88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1355_l1334_DUPLICATE_2c0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1350_l1337_DUPLICATE_8ec4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1350_l1337_DUPLICATE_8ec4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1350_l1327_l1337_l1334_DUPLICATE_7265_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1345_c30_bd88_return_output;
     -- CAST_TO_uint8_t[uxn_opcodes_h_l1353_c21_ff03] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1353_c21_ff03_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l1353_c31_f4c2_return_output);

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c7_a636] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l1339_c3_8499] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_x <= VAR_CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output := CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1350_c7_6af6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1342_c3_f5e1] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_left;
     BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output := BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1350_c7_6af6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c7_a636] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_left := VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1342_c3_f5e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1353_c21_ff03_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l1339_c3_8499_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c7_a636_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c7_a636_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l1343_c11_3ebf] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output;

     -- t16_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1350_c7_6af6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1350_c7_6af6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1350_c7_6af6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- Submodule level 3
     VAR_tmp16_uxn_opcodes_h_l1343_c3_1378 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1343_c11_3ebf_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1350_c7_6af6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := VAR_tmp16_uxn_opcodes_h_l1343_c3_1378;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1348_c21_f3c2] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1348_c21_f3c2_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_tmp16_uxn_opcodes_h_l1343_c3_1378);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- t16_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- Submodule level 4
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1348_c21_f3c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1341_c7_d4b7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- t16_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1341_c7_d4b7_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- t16_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     t16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     t16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1337_c7_15c1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1337_c7_15c1_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1334_c7_e39f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- Submodule level 7
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_e39f_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1327_c2_a117] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output := result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1323_l1360_DUPLICATE_ca38 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1323_l1360_DUPLICATE_ca38_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c2_a117_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c2_a117_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1323_l1360_DUPLICATE_ca38_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1323_l1360_DUPLICATE_ca38_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
