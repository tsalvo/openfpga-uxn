-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 56
entity swp_0CLK_bf6dd460 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_bf6dd460;
architecture arch of swp_0CLK_bf6dd460 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2715_c6_ed8c]
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2715_c1_56b3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2715_c2_c2e8]
signal n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2716_c3_3295[uxn_opcodes_h_l2716_c3_3295]
signal printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2720_c11_1d76]
signal BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal t8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2720_c7_bd08]
signal n8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2723_c11_ec54]
signal BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2723_c7_e057]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2723_c7_e057]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2723_c7_e057]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2723_c7_e057]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2723_c7_e057]
signal result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2723_c7_e057]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2723_c7_e057]
signal t8_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2723_c7_e057]
signal n8_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2727_c11_d91a]
signal BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2727_c7_217f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2727_c7_217f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2727_c7_217f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2727_c7_217f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2727_c7_217f]
signal result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2727_c7_217f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2727_c7_217f]
signal n8_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2730_c11_013a]
signal BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2730_c7_b2e7]
signal n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2733_c30_3fbb]
signal sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_6ae7]
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2738_c7_5980]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2738_c7_5980]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_5980]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_5980]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2738_c7_5980]
signal result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2743_c11_99b7]
signal BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2743_c7_a26b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2743_c7_a26b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c
BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_left,
BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_right,
BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8
result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- t8_MUX_uxn_opcodes_h_l2715_c2_c2e8
t8_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- n8_MUX_uxn_opcodes_h_l2715_c2_c2e8
n8_MUX_uxn_opcodes_h_l2715_c2_c2e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond,
n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue,
n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse,
n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

-- printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295
printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295 : entity work.printf_uxn_opcodes_h_l2716_c3_3295_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_left,
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_right,
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08
result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- t8_MUX_uxn_opcodes_h_l2720_c7_bd08
t8_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- n8_MUX_uxn_opcodes_h_l2720_c7_bd08
n8_MUX_uxn_opcodes_h_l2720_c7_bd08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond,
n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue,
n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse,
n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54
BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_left,
BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_right,
BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057
result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057
result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057
result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057
result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057
result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- t8_MUX_uxn_opcodes_h_l2723_c7_e057
t8_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
t8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
t8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- n8_MUX_uxn_opcodes_h_l2723_c7_e057
n8_MUX_uxn_opcodes_h_l2723_c7_e057 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2723_c7_e057_cond,
n8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue,
n8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse,
n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a
BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_left,
BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_right,
BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f
result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f
result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f
result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f
result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- n8_MUX_uxn_opcodes_h_l2727_c7_217f
n8_MUX_uxn_opcodes_h_l2727_c7_217f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2727_c7_217f_cond,
n8_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue,
n8_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse,
n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a
BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_left,
BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_right,
BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7
result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7
result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7
result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7
result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- n8_MUX_uxn_opcodes_h_l2730_c7_b2e7
n8_MUX_uxn_opcodes_h_l2730_c7_b2e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond,
n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue,
n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse,
n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb
sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_ins,
sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_x,
sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_y,
sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_left,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_right,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980
result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_cond,
result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7
BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_left,
BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_right,
BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b
result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b
result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output,
 sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2717_c3_7fd7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2721_c3_403e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2725_c3_741d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2728_c3_e513 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_4bb9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2740_c3_db3b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2738_c7_5980_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2748_l2711_DUPLICATE_01f1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2721_c3_403e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2721_c3_403e;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_4bb9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_4bb9;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2717_c3_7fd7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2717_c3_7fd7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2728_c3_e513 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2728_c3_e513;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2740_c3_db3b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2740_c3_db3b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2725_c3_741d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2725_c3_741d;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2738_c7_5980] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2738_c7_5980_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_6ae7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2727_c11_d91a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2733_c30_3fbb] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_ins;
     sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_x;
     sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output := sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2730_c11_013a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2723_c11_ec54] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_left;
     BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output := BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2743_c11_99b7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2720_c11_1d76] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_left;
     BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output := BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2715_c6_ed8c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c6_ed8c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_1d76_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2723_c11_ec54_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2727_c11_d91a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2730_c11_013a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_6ae7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2743_c11_99b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2720_l2715_l2730_l2727_l2723_DUPLICATE_38c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2720_l2743_l2738_l2730_l2727_l2723_DUPLICATE_5d8c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_deaf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2720_l2715_l2743_l2738_l2727_l2723_DUPLICATE_ab93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2720_l2715_l2738_l2727_l2723_DUPLICATE_aa86_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2738_c7_5980_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2733_c30_3fbb_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2715_c1_56b3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output;

     -- t8_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     t8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     t8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- n8_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2738_c7_5980] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output := result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2738_c7_5980] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2743_c7_a26b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2743_c7_a26b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2738_c7_5980] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2715_c1_56b3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2743_c7_a26b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_5980] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;

     -- t8_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- printf_uxn_opcodes_h_l2716_c3_3295[uxn_opcodes_h_l2716_c3_3295] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2716_c3_3295_uxn_opcodes_h_l2716_c3_3295_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     n8_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     n8_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_5980] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_5980_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     -- t8_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2730_c7_b2e7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     n8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     n8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2730_c7_b2e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;
     -- n8_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2727_c7_217f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2727_c7_217f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- n8_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2723_c7_e057] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2723_c7_e057_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2720_c7_bd08] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_bd08_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2715_c2_c2e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2748_l2711_DUPLICATE_01f1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2748_l2711_DUPLICATE_01f1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c2_c2e8_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2748_l2711_DUPLICATE_01f1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2748_l2711_DUPLICATE_01f1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
