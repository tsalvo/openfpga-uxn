-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldr_0CLK_5cd52163 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_5cd52163;
architecture arch of ldr_0CLK_5cd52163 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1604_c6_4688]
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l1604_c2_fb81]
signal t8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1617_c11_52ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1617_c7_a350]
signal tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1617_c7_a350]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1617_c7_a350]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1617_c7_a350]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1617_c7_a350]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1617_c7_a350]
signal result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1617_c7_a350]
signal result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l1617_c7_a350]
signal t8_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1620_c11_324d]
signal BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l1620_c7_8c40]
signal t8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1622_c30_ea46]
signal sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output : signed(3 downto 0);

-- u16_add_u8_as_i8[uxn_opcodes_h_l1623_c22_85a9]
signal u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u16 : unsigned(15 downto 0);
signal u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u8 : unsigned(7 downto 0);
signal u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1625_c11_9e7e]
signal BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1625_c7_7664]
signal tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1625_c7_7664]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1625_c7_7664]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1625_c7_7664]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1625_c7_7664]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1625_c7_7664]
signal result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1628_c11_c671]
signal BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1628_c7_efb7]
signal tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1628_c7_efb7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1628_c7_efb7]
signal result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1628_c7_efb7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1628_c7_efb7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_ram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.u16_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_left,
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_right,
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81
tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81
result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81
result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81
result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- t8_MUX_uxn_opcodes_h_l1604_c2_fb81
t8_MUX_uxn_opcodes_h_l1604_c2_fb81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond,
t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue,
t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse,
t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed
BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1617_c7_a350
tmp8_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350
result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350
result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350
result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350
result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350
result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- t8_MUX_uxn_opcodes_h_l1617_c7_a350
t8_MUX_uxn_opcodes_h_l1617_c7_a350 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1617_c7_a350_cond,
t8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue,
t8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse,
t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_left,
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_right,
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40
tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40
result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- t8_MUX_uxn_opcodes_h_l1620_c7_8c40
t8_MUX_uxn_opcodes_h_l1620_c7_8c40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond,
t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue,
t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse,
t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46
sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_ins,
sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_x,
sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_y,
sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output);

-- u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9
u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9 : entity work.u16_add_u8_as_i8_0CLK_e595f783 port map (
u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u16,
u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u8,
u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e
BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_left,
BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_right,
BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1625_c7_7664
tmp8_MUX_uxn_opcodes_h_l1625_c7_7664 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_cond,
tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue,
tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse,
tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664
result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664
result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664
result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664
result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_cond,
result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671
BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_left,
BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_right,
BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7
tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_cond,
tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue,
tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse,
tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7
result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7
result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7
result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output,
 tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output,
 tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output,
 tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output,
 sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output,
 u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output,
 tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output,
 tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_b402 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1609_c3_15c6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1618_c3_82f1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output : signed(3 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u16 : unsigned(15 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u8 : unsigned(7 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1626_c3_e719 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1631_c3_1847 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1617_l1620_l1604_DUPLICATE_9022_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1625_l1617_DUPLICATE_d239_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1625_l1628_l1620_DUPLICATE_1312_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1600_l1636_DUPLICATE_cec8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_b402 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_b402;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1631_c3_1847 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1631_c3_1847;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1626_c3_e719 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1626_c3_e719;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1609_c3_15c6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1609_c3_15c6;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1618_c3_82f1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1618_c3_82f1;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_ins := VAR_ins;
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u16 := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_previous_stack_read;
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u8 := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1617_c11_52ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1625_l1628_l1620_DUPLICATE_1312 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1625_l1628_l1620_DUPLICATE_1312_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1617_l1620_l1604_DUPLICATE_9022 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1617_l1620_l1604_DUPLICATE_9022_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l1622_c30_ea46] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_ins;
     sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_x;
     sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output := sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1604_c6_4688] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_left;
     BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output := BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;

     -- u16_add_u8_as_i8[uxn_opcodes_h_l1623_c22_85a9] LATENCY=0
     -- Inputs
     u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u16 <= VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u16;
     u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u8 <= VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_u8;
     -- Outputs
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output := u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1620_c11_324d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1625_c11_9e7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1628_c11_c671] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_left;
     BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output := BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1625_l1617_DUPLICATE_d239 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1625_l1617_DUPLICATE_d239_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_4688_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1617_c11_52ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_324d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1625_c11_9e7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1628_c11_c671_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1625_l1617_DUPLICATE_d239_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1625_l1617_DUPLICATE_d239_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1617_l1620_l1604_DUPLICATE_9022_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1617_l1620_l1604_DUPLICATE_9022_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1617_l1620_l1604_DUPLICATE_9022_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_1b07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1625_l1617_l1628_l1620_DUPLICATE_bb97_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1625_l1628_l1620_DUPLICATE_1312_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1625_l1628_l1620_DUPLICATE_1312_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1625_l1628_l1620_DUPLICATE_1312_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1625_l1620_l1617_l1604_l1628_DUPLICATE_3cfb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1604_c2_fb81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1622_c30_ea46_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue := VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1623_c22_85a9_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1628_c7_efb7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1628_c7_efb7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1625_c7_7664] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1628_c7_efb7] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_cond;
     tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output := tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1628_c7_efb7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1628_c7_efb7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- t8_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1628_c7_efb7_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1625_c7_7664] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1625_c7_7664] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1625_c7_7664] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output := result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1625_c7_7664] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_cond;
     tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output := tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1625_c7_7664] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;

     -- t8_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     t8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     t8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1625_c7_7664_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- t8_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1620_c7_8c40] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_8c40_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1617_c7_a350] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1617_c7_a350_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1604_c2_fb81] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1600_l1636_DUPLICATE_cec8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1600_l1636_DUPLICATE_cec8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_fb81_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1600_l1636_DUPLICATE_cec8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1600_l1636_DUPLICATE_cec8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
