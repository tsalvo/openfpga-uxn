-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity ldr_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_f74745d5;
architecture arch of ldr_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1600_c6_e094]
signal BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1600_c2_1caa]
signal t8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1613_c11_0225]
signal BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1613_c7_827b]
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1613_c7_827b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1613_c7_827b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1613_c7_827b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1613_c7_827b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1613_c7_827b]
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1613_c7_827b]
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1613_c7_827b]
signal t8_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1616_c11_a356]
signal BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1616_c7_ca9c]
signal t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1618_c30_a015]
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1619_c22_ff98]
signal BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1621_c11_e078]
signal BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1621_c7_d153]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1621_c7_d153]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1621_c7_d153]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1621_c7_d153]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1621_c7_d153]
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1621_c7_d153]
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1624_c11_21a8]
signal BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1624_c7_967c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1624_c7_967c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1624_c7_967c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1624_c7_967c]
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1624_c7_967c]
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(7 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a906( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.u8_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_left,
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_right,
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa
tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- t8_MUX_uxn_opcodes_h_l1600_c2_1caa
t8_MUX_uxn_opcodes_h_l1600_c2_1caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond,
t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue,
t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse,
t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_left,
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_right,
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1613_c7_827b
tmp8_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- t8_MUX_uxn_opcodes_h_l1613_c7_827b
t8_MUX_uxn_opcodes_h_l1613_c7_827b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1613_c7_827b_cond,
t8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue,
t8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse,
t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_left,
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_right,
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c
tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- t8_MUX_uxn_opcodes_h_l1616_c7_ca9c
t8_MUX_uxn_opcodes_h_l1616_c7_ca9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond,
t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue,
t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse,
t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1618_c30_a015
sp_relative_shift_uxn_opcodes_h_l1618_c30_a015 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_ins,
sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_x,
sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_y,
sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_left,
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_right,
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_left,
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_right,
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_cond,
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1621_c7_d153
tmp8_MUX_uxn_opcodes_h_l1621_c7_d153 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_cond,
tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue,
tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse,
tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_left,
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_right,
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1624_c7_967c
tmp8_MUX_uxn_opcodes_h_l1624_c7_967c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_cond,
tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output,
 tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_40bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1605_c3_473d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_816d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1619_c3_c5cc : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1619_c27_d5bd_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1622_c3_4202 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1627_c3_ad7b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_3c24_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_114a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_8e1b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1596_l1632_DUPLICATE_665a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_40bb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_40bb;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1605_c3_473d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1605_c3_473d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_816d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_816d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1622_c3_4202 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1622_c3_4202;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1627_c3_ad7b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1627_c3_ad7b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1613_c11_0225] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_left;
     BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output := BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1618_c30_a015] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_ins;
     sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_x;
     sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output := sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_8e1b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_8e1b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1616_c11_a356] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_left;
     BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output := BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_114a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_114a_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_3c24 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_3c24_return_output := result.u16_value;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1619_c27_d5bd] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1619_c27_d5bd_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1600_c6_e094] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_left;
     BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output := BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1621_c11_e078] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_left;
     BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output := BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1624_c11_21a8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_e094_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0225_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_a356_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_e078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_21a8_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1619_c27_d5bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_114a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_114a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_3c24_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_3c24_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_3c24_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_cc89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_145e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_8e1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_8e1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_8e1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1624_l1621_l1616_l1613_l1600_DUPLICATE_73eb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1600_c2_1caa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_a015_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1624_c7_967c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_cond;
     tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output := tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1621_c7_d153] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1624_c7_967c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1624_c7_967c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1619_c22_ff98] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1624_c7_967c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1624_c7_967c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1619_c3_c5cc := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_ff98_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_967c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1619_c3_c5cc;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1621_c7_d153] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1621_c7_d153] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output := result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1621_c7_d153] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1621_c7_d153] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;

     -- t8_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     t8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     t8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1621_c7_d153] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_cond;
     tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output := tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_d153_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1616_c7_ca9c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_ca9c_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1613_c7_827b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_827b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1600_c2_1caa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1596_l1632_DUPLICATE_665a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1596_l1632_DUPLICATE_665a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a906(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_1caa_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1596_l1632_DUPLICATE_665a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1596_l1632_DUPLICATE_665a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
