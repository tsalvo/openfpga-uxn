-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity add_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end add_0CLK_bacf6a1d;
architecture arch of add_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l790_c6_fe02]
signal BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l790_c1_ed4a]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal n8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal t8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l790_c2_b0e8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l791_c3_33a6[uxn_opcodes_h_l791_c3_33a6]
signal printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l795_c11_c3b2]
signal BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal n8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal t8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l795_c7_d8e8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l798_c11_84e7]
signal BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l798_c7_5268]
signal n8_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l798_c7_5268]
signal t8_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l798_c7_5268]
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l798_c7_5268]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l798_c7_5268]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l798_c7_5268]
signal result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l798_c7_5268]
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l798_c7_5268]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l801_c11_aa67]
signal BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l801_c7_82ed]
signal n8_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l801_c7_82ed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l801_c7_82ed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l801_c7_82ed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l801_c7_82ed]
signal result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l801_c7_82ed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l801_c7_82ed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l804_c30_4d6d]
signal sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l807_c21_1cc5]
signal BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l809_c11_69e2]
signal BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l809_c7_82ba]
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l809_c7_82ba]
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l809_c7_82ba]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02
BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_left,
BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_right,
BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output);

-- n8_MUX_uxn_opcodes_h_l790_c2_b0e8
n8_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- t8_MUX_uxn_opcodes_h_l790_c2_b0e8
t8_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8
result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8
result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8
result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8
result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

-- printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6
printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6 : entity work.printf_uxn_opcodes_h_l791_c3_33a6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2
BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_left,
BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_right,
BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output);

-- n8_MUX_uxn_opcodes_h_l795_c7_d8e8
n8_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- t8_MUX_uxn_opcodes_h_l795_c7_d8e8
t8_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8
result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8
result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7
BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_left,
BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_right,
BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output);

-- n8_MUX_uxn_opcodes_h_l798_c7_5268
n8_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l798_c7_5268_cond,
n8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
n8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- t8_MUX_uxn_opcodes_h_l798_c7_5268
t8_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l798_c7_5268_cond,
t8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
t8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268
result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268
result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_cond,
result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268
result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67
BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_left,
BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_right,
BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output);

-- n8_MUX_uxn_opcodes_h_l801_c7_82ed
n8_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
n8_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
n8_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed
result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed
result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed
result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed
result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed
result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output);

-- sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d
sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_ins,
sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_x,
sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_y,
sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5
BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5 : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_left,
BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_right,
BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2
BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_left,
BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_right,
BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output,
 n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output,
 n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output,
 n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output,
 n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output,
 sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l792_c3_cb18 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l796_c3_dde4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l806_c3_e79a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l807_c3_62c7 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l798_l801_DUPLICATE_06a9_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l815_l786_DUPLICATE_3ec8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l792_c3_cb18 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l792_c3_cb18;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l806_c3_e79a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l806_c3_e79a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l796_c3_dde4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l796_c3_dde4;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l798_l801_DUPLICATE_06a9 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l798_l801_DUPLICATE_06a9_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l804_c30_4d6d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_ins;
     sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_x;
     sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output := sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l798_c11_84e7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_left;
     BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output := BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l795_c11_c3b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l790_c6_fe02] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_left;
     BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output := BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l809_c11_69e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l801_c11_aa67] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_left;
     BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output := BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41_return_output := result.is_opc_done;

     -- BIN_OP_PLUS[uxn_opcodes_h_l807_c21_1cc5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_left;
     BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output := BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c6_fe02_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_c3b2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c11_84e7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l801_c11_aa67_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_69e2_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l807_c3_62c7 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l807_c21_1cc5_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_e143_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l795_l809_l798_l801_DUPLICATE_ab41_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_dc8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l795_l809_l798_l790_DUPLICATE_a8b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l798_l801_DUPLICATE_06a9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l798_l801_DUPLICATE_06a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l795_l798_l790_l801_DUPLICATE_1ed9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l804_c30_4d6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue := VAR_result_u8_value_uxn_opcodes_h_l807_c3_62c7;
     -- t8_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     t8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     t8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output := t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l809_c7_82ba] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- n8_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     n8_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     n8_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l809_c7_82ba] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l809_c7_82ba] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l790_c1_ed4a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l790_c1_ed4a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_n8_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_82ba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_82ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_82ba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output := result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- printf_uxn_opcodes_h_l791_c3_33a6[uxn_opcodes_h_l791_c3_33a6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l791_c3_33a6_uxn_opcodes_h_l791_c3_33a6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- t8_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l801_c7_82ed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;

     -- n8_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     n8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     n8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output := n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l801_c7_82ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- t8_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- n8_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l798_c7_5268] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c7_5268_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l795_c7_d8e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- n8_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_d8e8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l790_c2_b0e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l815_l786_DUPLICATE_3ec8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l815_l786_DUPLICATE_3ec8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l790_c2_b0e8_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l815_l786_DUPLICATE_3ec8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l815_l786_DUPLICATE_3ec8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
