-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity inc_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_66ba3dc0;
architecture arch of inc_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1489_c6_463f]
signal BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1489_c1_5f1c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1489_c2_a4eb]
signal t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1490_c3_9231[uxn_opcodes_h_l1490_c3_9231]
signal printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1495_c11_4244]
signal BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1495_c7_03ff]
signal t8_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1498_c11_78bd]
signal BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1498_c7_a13a]
signal t8_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1502_c32_26df]
signal BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1502_c32_405d]
signal BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1502_c32_ba14]
signal MUX_uxn_opcodes_h_l1502_c32_ba14_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1502_c32_ba14_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1502_c32_ba14_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1502_c32_ba14_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1504_c11_3d79]
signal BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1504_c7_ea22]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1504_c7_ea22]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1504_c7_ea22]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1504_c7_ea22]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1504_c7_ea22]
signal result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1508_c24_8a0c]
signal BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1510_c11_645b]
signal BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1510_c7_2e05]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1510_c7_2e05]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_1ade( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.is_stack_read := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.stack_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f
BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_left,
BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_right,
BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb
result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- t8_MUX_uxn_opcodes_h_l1489_c2_a4eb
t8_MUX_uxn_opcodes_h_l1489_c2_a4eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond,
t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue,
t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse,
t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

-- printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231
printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231 : entity work.printf_uxn_opcodes_h_l1490_c3_9231_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244
BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_left,
BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_right,
BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff
result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff
result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff
result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff
result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff
result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- t8_MUX_uxn_opcodes_h_l1495_c7_03ff
t8_MUX_uxn_opcodes_h_l1495_c7_03ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1495_c7_03ff_cond,
t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue,
t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse,
t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd
BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_left,
BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_right,
BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a
result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a
result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a
result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a
result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a
result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- t8_MUX_uxn_opcodes_h_l1498_c7_a13a
t8_MUX_uxn_opcodes_h_l1498_c7_a13a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1498_c7_a13a_cond,
t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue,
t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse,
t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df
BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_left,
BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_right,
BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d
BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_left,
BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_right,
BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output);

-- MUX_uxn_opcodes_h_l1502_c32_ba14
MUX_uxn_opcodes_h_l1502_c32_ba14 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1502_c32_ba14_cond,
MUX_uxn_opcodes_h_l1502_c32_ba14_iftrue,
MUX_uxn_opcodes_h_l1502_c32_ba14_iffalse,
MUX_uxn_opcodes_h_l1502_c32_ba14_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79
BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_left,
BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_right,
BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22
result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22
result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22
result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22
result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_cond,
result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c
BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_left,
BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_right,
BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b
BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_left,
BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_right,
BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05
result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05
result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output,
 MUX_uxn_opcodes_h_l1502_c32_ba14_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1492_c3_fe57 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1496_c3_f63b : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1507_c3_b80a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1508_c3_1d9e : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1489_l1504_l1495_DUPLICATE_65e6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1498_l1489_l1495_DUPLICATE_40b1_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1498_l1495_DUPLICATE_976d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1498_l1504_DUPLICATE_8a6a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l1515_l1485_DUPLICATE_bbf8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1492_c3_fe57 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1492_c3_fe57;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_right := to_unsigned(128, 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1507_c3_b80a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1507_c3_b80a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1496_c3_f63b := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1496_c3_f63b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_right := to_unsigned(3, 2);
     VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := t8;
     -- BIN_OP_PLUS[uxn_opcodes_h_l1508_c24_8a0c] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1498_l1495_DUPLICATE_976d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1498_l1495_DUPLICATE_976d_return_output := result.is_stack_read;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1495_c11_4244] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_left;
     BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output := BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1498_l1489_l1495_DUPLICATE_40b1 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1498_l1489_l1495_DUPLICATE_40b1_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1498_c11_78bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1498_l1504_DUPLICATE_8a6a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1498_l1504_DUPLICATE_8a6a_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1489_c6_463f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l1502_c32_26df] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_left;
     BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output := BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1510_c11_645b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1489_l1504_l1495_DUPLICATE_65e6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1489_l1504_l1495_DUPLICATE_65e6_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1504_c11_3d79] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_left;
     BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output := BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1502_c32_26df_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c6_463f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1495_c11_4244_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1498_c11_78bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1504_c11_3d79_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1510_c11_645b_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1508_c3_1d9e := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1508_c24_8a0c_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1498_l1489_l1495_DUPLICATE_40b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1498_l1489_l1495_DUPLICATE_40b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1498_l1489_l1495_DUPLICATE_40b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1498_l1504_l1495_l1510_DUPLICATE_7d89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1489_l1504_l1495_DUPLICATE_65e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1489_l1504_l1495_DUPLICATE_65e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1489_l1504_l1495_DUPLICATE_65e6_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1498_l1495_DUPLICATE_976d_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1498_l1495_DUPLICATE_976d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1498_l1489_l1495_l1510_DUPLICATE_17f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1498_l1504_DUPLICATE_8a6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1498_l1504_DUPLICATE_8a6a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1498_l1489_l1504_l1495_DUPLICATE_9a2e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1508_c3_1d9e;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1504_c7_ea22] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1504_c7_ea22] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1489_c1_5f1c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1504_c7_ea22] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output := result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1502_c32_405d] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_left;
     BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output := BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1510_c7_2e05] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1510_c7_2e05] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1502_c32_405d_return_output;
     VAR_printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1489_c1_5f1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1510_c7_2e05_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- t8_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- printf_uxn_opcodes_h_l1490_c3_9231[uxn_opcodes_h_l1490_c3_9231] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1490_c3_9231_uxn_opcodes_h_l1490_c3_9231_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1504_c7_ea22] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;

     -- MUX[uxn_opcodes_h_l1502_c32_ba14] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1502_c32_ba14_cond <= VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_cond;
     MUX_uxn_opcodes_h_l1502_c32_ba14_iftrue <= VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_iftrue;
     MUX_uxn_opcodes_h_l1502_c32_ba14_iffalse <= VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_return_output := MUX_uxn_opcodes_h_l1502_c32_ba14_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1504_c7_ea22] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue := VAR_MUX_uxn_opcodes_h_l1502_c32_ba14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1504_c7_ea22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- t8_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1498_c7_a13a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1498_c7_a13a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1495_c7_03ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1495_c7_03ff_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1489_c2_a4eb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l1515_l1485_DUPLICATE_bbf8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l1515_l1485_DUPLICATE_bbf8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1ade(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1489_c2_a4eb_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l1515_l1485_DUPLICATE_bbf8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l1515_l1485_DUPLICATE_bbf8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
