-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity add2_0CLK_06b39b76 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end add2_0CLK_06b39b76;
architecture arch of add2_0CLK_06b39b76 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l814_c6_4728]
signal BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l814_c2_efa7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l814_c2_efa7]
signal n16_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l814_c2_efa7]
signal tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l814_c2_efa7]
signal t16_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l822_c11_dfcf]
signal BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal n16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l822_c7_1e5a]
signal t16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l825_c11_1b37]
signal BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l825_c7_201e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l825_c7_201e]
signal n16_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l825_c7_201e]
signal tmp16_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l825_c7_201e]
signal t16_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l828_c30_8086]
signal sp_relative_shift_uxn_opcodes_h_l828_c30_8086_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l828_c30_8086_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l828_c30_8086_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l830_c11_2c56]
signal BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l830_c7_66eb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l830_c7_66eb]
signal result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l830_c7_66eb]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l830_c7_66eb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l830_c7_66eb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l830_c7_66eb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l830_c7_66eb]
signal n16_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l830_c7_66eb]
signal tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l832_c11_6523]
signal BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_right : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l838_c11_4fe5]
signal BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l838_c7_01ea]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l838_c7_01ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l838_c7_01ea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728
BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_left,
BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_right,
BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7
result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7
result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7
result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7
result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7
result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- n16_MUX_uxn_opcodes_h_l814_c2_efa7
n16_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
n16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
n16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- tmp16_MUX_uxn_opcodes_h_l814_c2_efa7
tmp16_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- t16_MUX_uxn_opcodes_h_l814_c2_efa7
t16_MUX_uxn_opcodes_h_l814_c2_efa7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l814_c2_efa7_cond,
t16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue,
t16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse,
t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf
BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_left,
BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_right,
BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a
result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a
result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a
result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a
result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a
result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- n16_MUX_uxn_opcodes_h_l822_c7_1e5a
n16_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a
tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- t16_MUX_uxn_opcodes_h_l822_c7_1e5a
t16_MUX_uxn_opcodes_h_l822_c7_1e5a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond,
t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue,
t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse,
t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37
BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_left,
BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_right,
BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e
result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e
result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e
result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e
result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e
result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- n16_MUX_uxn_opcodes_h_l825_c7_201e
n16_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l825_c7_201e_cond,
n16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
n16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- tmp16_MUX_uxn_opcodes_h_l825_c7_201e
tmp16_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l825_c7_201e_cond,
tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- t16_MUX_uxn_opcodes_h_l825_c7_201e
t16_MUX_uxn_opcodes_h_l825_c7_201e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l825_c7_201e_cond,
t16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue,
t16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse,
t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l828_c30_8086
sp_relative_shift_uxn_opcodes_h_l828_c30_8086 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l828_c30_8086_ins,
sp_relative_shift_uxn_opcodes_h_l828_c30_8086_x,
sp_relative_shift_uxn_opcodes_h_l828_c30_8086_y,
sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56
BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_left,
BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_right,
BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb
result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb
result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb
result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb
result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- n16_MUX_uxn_opcodes_h_l830_c7_66eb
n16_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
n16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
n16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- tmp16_MUX_uxn_opcodes_h_l830_c7_66eb
tmp16_MUX_uxn_opcodes_h_l830_c7_66eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_cond,
tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue,
tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse,
tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523
BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523 : entity work.BIN_OP_PLUS_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_left,
BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_right,
BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5
BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_left,
BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_right,
BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea
result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea
result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output,
 sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l819_c3_948d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l823_c3_ed3d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l835_c3_22e7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_uxn_opcodes_h_l832_c3_51b5 : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l822_l830_l814_DUPLICATE_8162_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l825_l822_l814_DUPLICATE_ff81_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l825_l830_DUPLICATE_cc73_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l844_l810_DUPLICATE_1379_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l835_c3_22e7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l835_c3_22e7;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_right := to_unsigned(4, 3);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l819_c3_948d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l819_c3_948d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l823_c3_ed3d := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l823_c3_ed3d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := t16;
     VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := tmp16;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l825_l830_DUPLICATE_cc73 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l825_l830_DUPLICATE_cc73_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l838_c11_4fe5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_left;
     BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output := BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l825_c11_1b37] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_left;
     BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output := BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l822_l830_l814_DUPLICATE_8162 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l822_l830_l814_DUPLICATE_8162_return_output := result.is_sp_shift;

     -- BIN_OP_PLUS[uxn_opcodes_h_l832_c11_6523] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_left;
     BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output := BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e_return_output := result.u16_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l825_l822_l814_DUPLICATE_ff81 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l825_l822_l814_DUPLICATE_ff81_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l830_c11_2c56] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_left;
     BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output := BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_EQ[uxn_opcodes_h_l822_c11_dfcf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_left;
     BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output := BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l814_c6_4728] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_left;
     BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output := BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l828_c30_8086] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l828_c30_8086_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_ins;
     sp_relative_shift_uxn_opcodes_h_l828_c30_8086_x <= VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_x;
     sp_relative_shift_uxn_opcodes_h_l828_c30_8086_y <= VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output := sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l814_c6_4728_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l822_c11_dfcf_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l825_c11_1b37_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l830_c11_2c56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l838_c11_4fe5_return_output;
     VAR_tmp16_uxn_opcodes_h_l832_c3_51b5 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l832_c11_6523_return_output, 16);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l825_l822_l814_DUPLICATE_ff81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l825_l822_l814_DUPLICATE_ff81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l825_l822_l814_DUPLICATE_ff81_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l825_l822_l830_l814_DUPLICATE_302e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_bacc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l822_l830_l814_DUPLICATE_8162_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l822_l830_l814_DUPLICATE_8162_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l822_l830_l814_DUPLICATE_8162_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l825_l822_l830_l838_DUPLICATE_184b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l825_l822_l838_l814_DUPLICATE_3a55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l825_l830_DUPLICATE_cc73_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l825_l830_DUPLICATE_cc73_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l828_c30_8086_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := VAR_tmp16_uxn_opcodes_h_l832_c3_51b5;
     VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue := VAR_tmp16_uxn_opcodes_h_l832_c3_51b5;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l838_c7_01ea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l838_c7_01ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output;

     -- n16_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     n16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     n16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l838_c7_01ea] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- t16_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     t16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     t16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output := t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_n16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l838_c7_01ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l838_c7_01ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l838_c7_01ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- t16_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- n16_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     n16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     n16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output := n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output := tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l830_c7_66eb] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_n16_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l830_c7_66eb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_t16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     -- t16_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     t16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     t16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- n16_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l825_c7_201e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_n16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l825_c7_201e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- n16_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     n16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     n16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l822_c7_1e5a] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l822_c7_1e5a_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l814_c2_efa7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l844_l810_DUPLICATE_1379 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l844_l810_DUPLICATE_1379_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l814_c2_efa7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l814_c2_efa7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l844_l810_DUPLICATE_1379_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l844_l810_DUPLICATE_1379_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
