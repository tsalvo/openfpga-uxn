-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1185_c6_f8d8]
signal BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1185_c2_3468]
signal t8_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1185_c2_3468]
signal n8_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1185_c2_3468]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1198_c11_4f73]
signal BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1198_c7_e6ec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1201_c11_b69d]
signal BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal t8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal n8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1201_c7_3f15]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1204_c11_fd86]
signal BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1204_c7_950e]
signal n8_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1204_c7_950e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1204_c7_950e]
signal result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1204_c7_950e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1204_c7_950e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1204_c7_950e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1206_c30_94af]
signal sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1209_c21_37ea]
signal BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1209_c21_7f64]
signal MUX_uxn_opcodes_h_l1209_c21_7f64_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1209_c21_7f64_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1209_c21_7f64_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1209_c21_7f64_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8
BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_left,
BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_right,
BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output);

-- t8_MUX_uxn_opcodes_h_l1185_c2_3468
t8_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
t8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
t8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- n8_MUX_uxn_opcodes_h_l1185_c2_3468
n8_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
n8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
n8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468
result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468
result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468
result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468
result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73
BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_left,
BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_right,
BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output);

-- t8_MUX_uxn_opcodes_h_l1198_c7_e6ec
t8_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- n8_MUX_uxn_opcodes_h_l1198_c7_e6ec
n8_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec
result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec
result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec
result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec
result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d
BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_left,
BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_right,
BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output);

-- t8_MUX_uxn_opcodes_h_l1201_c7_3f15
t8_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- n8_MUX_uxn_opcodes_h_l1201_c7_3f15
n8_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15
result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15
result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15
result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15
result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86
BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_left,
BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_right,
BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output);

-- n8_MUX_uxn_opcodes_h_l1204_c7_950e
n8_MUX_uxn_opcodes_h_l1204_c7_950e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1204_c7_950e_cond,
n8_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue,
n8_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse,
n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e
result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e
result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e
result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1206_c30_94af
sp_relative_shift_uxn_opcodes_h_l1206_c30_94af : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_ins,
sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_x,
sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_y,
sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea
BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_left,
BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_right,
BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output);

-- MUX_uxn_opcodes_h_l1209_c21_7f64
MUX_uxn_opcodes_h_l1209_c21_7f64 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1209_c21_7f64_cond,
MUX_uxn_opcodes_h_l1209_c21_7f64_iftrue,
MUX_uxn_opcodes_h_l1209_c21_7f64_iffalse,
MUX_uxn_opcodes_h_l1209_c21_7f64_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output,
 t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output,
 t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output,
 t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output,
 n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output,
 sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output,
 MUX_uxn_opcodes_h_l1209_c21_7f64_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1190_c3_1461 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1195_c3_b310 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1199_c3_18c8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1208_c3_8151 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_4f1c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_c9be_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_5ac4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1204_l1201_DUPLICATE_3596_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1213_l1181_DUPLICATE_f1a9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1190_c3_1461 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1190_c3_1461;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1199_c3_18c8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1199_c3_18c8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1195_c3_b310 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1195_c3_b310;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1208_c3_8151 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1208_c3_8151;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1204_c11_fd86] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_left;
     BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output := BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1185_c2_3468_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1206_c30_94af] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_ins;
     sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_x;
     sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output := sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_c9be LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_c9be_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1185_c6_f8d8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_5ac4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_5ac4_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_4f1c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_4f1c_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1185_c2_3468_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1185_c2_3468_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1209_c21_37ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1198_c11_4f73] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_left;
     BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output := BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1204_l1201_DUPLICATE_3596 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1204_l1201_DUPLICATE_3596_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1201_c11_b69d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1185_c2_3468_return_output := result.is_ram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c6_f8d8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1198_c11_4f73_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1201_c11_b69d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c11_fd86_return_output;
     VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1209_c21_37ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_c9be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_c9be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_c9be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_4f1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_4f1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_4f1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_5ac4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_5ac4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1204_l1198_l1201_DUPLICATE_5ac4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1204_l1201_DUPLICATE_3596_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1204_l1201_DUPLICATE_3596_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1204_l1198_l1201_DUPLICATE_9a5b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1185_c2_3468_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1185_c2_3468_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1185_c2_3468_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1185_c2_3468_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1206_c30_94af_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- MUX[uxn_opcodes_h_l1209_c21_7f64] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1209_c21_7f64_cond <= VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_cond;
     MUX_uxn_opcodes_h_l1209_c21_7f64_iftrue <= VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_iftrue;
     MUX_uxn_opcodes_h_l1209_c21_7f64_iffalse <= VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_return_output := MUX_uxn_opcodes_h_l1209_c21_7f64_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1204_c7_950e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1204_c7_950e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1204_c7_950e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1204_c7_950e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1204_c7_950e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1204_c7_950e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_cond;
     n8_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue;
     n8_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output := n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue := VAR_MUX_uxn_opcodes_h_l1209_c21_7f64_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1204_c7_950e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- t8_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- n8_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1204_c7_950e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- n8_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1201_c7_3f15] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output := result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;

     -- t8_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     t8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     t8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1201_c7_3f15_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;
     -- n8_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     n8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     n8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1198_c7_e6ec] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output := result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1198_c7_e6ec_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1185_c2_3468] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output := result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1213_l1181_DUPLICATE_f1a9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1213_l1181_DUPLICATE_f1a9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c2_3468_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1185_c2_3468_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1213_l1181_DUPLICATE_f1a9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1213_l1181_DUPLICATE_f1a9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
