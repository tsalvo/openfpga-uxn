-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_64d180f1;
architecture arch of eor_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1077_c6_8b60]
signal BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal n8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal t8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1077_c2_79a1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1090_c11_e6f9]
signal BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal n8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal t8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1090_c7_c96d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1093_c11_7a55]
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal n8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal t8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c7_c84c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1096_c11_f0dc]
signal BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1096_c7_b7a8]
signal n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1096_c7_b7a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1096_c7_b7a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1096_c7_b7a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1096_c7_b7a8]
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1096_c7_b7a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1098_c30_3bb5]
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1101_c21_61ea]
signal BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_left,
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_right,
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output);

-- n8_MUX_uxn_opcodes_h_l1077_c2_79a1
n8_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- t8_MUX_uxn_opcodes_h_l1077_c2_79a1
t8_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_left,
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_right,
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output);

-- n8_MUX_uxn_opcodes_h_l1090_c7_c96d
n8_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- t8_MUX_uxn_opcodes_h_l1090_c7_c96d
t8_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_left,
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_right,
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output);

-- n8_MUX_uxn_opcodes_h_l1093_c7_c84c
n8_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- t8_MUX_uxn_opcodes_h_l1093_c7_c84c
t8_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_left,
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_right,
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output);

-- n8_MUX_uxn_opcodes_h_l1096_c7_b7a8
n8_MUX_uxn_opcodes_h_l1096_c7_b7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond,
n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue,
n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse,
n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5
sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_ins,
sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_x,
sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_y,
sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_left,
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_right,
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output,
 n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output,
 n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output,
 n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output,
 n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output,
 sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1082_c3_df6e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1087_c3_cc61 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1091_c3_bd53 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1100_c3_59de : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_875a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_355f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_c074_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1093_l1096_DUPLICATE_8175_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1105_l1073_DUPLICATE_1aa2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1100_c3_59de := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1100_c3_59de;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_right := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1082_c3_df6e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1082_c3_df6e;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1087_c3_cc61 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1087_c3_cc61;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1091_c3_bd53 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1091_c3_bd53;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_875a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_875a_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output := result.is_ram_write;

     -- BIN_OP_XOR[uxn_opcodes_h_l1101_c21_61ea] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_left;
     BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output := BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1096_c11_f0dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_left;
     BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output := BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_355f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_355f_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1098_c30_3bb5] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_ins;
     sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_x;
     sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output := sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_c074 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_c074_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1077_c6_8b60] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_left;
     BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output := BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1090_c11_e6f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1093_c11_7a55] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_left;
     BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output := BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1093_l1096_DUPLICATE_8175 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1093_l1096_DUPLICATE_8175_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_8b60_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_e6f9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_7a55_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_f0dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_61ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_875a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_875a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_875a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_355f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_355f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_355f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_c074_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_c074_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1093_l1096_l1090_DUPLICATE_c074_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1093_l1096_DUPLICATE_8175_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1093_l1096_DUPLICATE_8175_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1093_l1077_l1096_l1090_DUPLICATE_e019_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1077_c2_79a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_3bb5_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1096_c7_b7a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1096_c7_b7a8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond <= VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond;
     n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue;
     n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output := n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1096_c7_b7a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1096_c7_b7a8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1096_c7_b7a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1096_c7_b7a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_b7a8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c7_c84c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_c84c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- n8_MUX[uxn_opcodes_h_l1090_c7_c96d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_cond;
     n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iftrue;
     n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output := n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_c96d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1077_c2_79a1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_cond;
     n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iftrue;
     n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output := n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1105_l1073_DUPLICATE_1aa2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1105_l1073_DUPLICATE_1aa2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_79a1_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1105_l1073_DUPLICATE_1aa2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1105_l1073_DUPLICATE_1aa2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
