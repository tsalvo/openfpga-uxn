-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 34
entity sth_0CLK_02ab8d09 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_02ab8d09;
architecture arch of sth_0CLK_02ab8d09 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2146_c6_de3d]
signal BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2146_c2_ee74]
signal t8_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2153_c11_adc8]
signal BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2153_c7_55d2]
signal t8_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2156_c30_9b72]
signal sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2158_c11_2195]
signal BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2158_c7_f092]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2158_c7_f092]
signal t8_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2166_c11_c6d2]
signal BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2166_c7_a66e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2166_c7_a66e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2166_c7_a66e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2166_c7_a66e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5c64( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d
BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_left,
BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_right,
BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74
result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74
result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74
result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74
result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74
result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- t8_MUX_uxn_opcodes_h_l2146_c2_ee74
t8_MUX_uxn_opcodes_h_l2146_c2_ee74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2146_c2_ee74_cond,
t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue,
t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse,
t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8
BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_left,
BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_right,
BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2
result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2
result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2
result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2
result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- t8_MUX_uxn_opcodes_h_l2153_c7_55d2
t8_MUX_uxn_opcodes_h_l2153_c7_55d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2153_c7_55d2_cond,
t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue,
t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse,
t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72
sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_ins,
sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_x,
sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_y,
sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195
BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_left,
BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_right,
BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092
result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092
result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092
result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092
result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092
result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- t8_MUX_uxn_opcodes_h_l2158_c7_f092
t8_MUX_uxn_opcodes_h_l2158_c7_f092 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2158_c7_f092_cond,
t8_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue,
t8_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse,
t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2
BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_left,
BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_right,
BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e
result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e
result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e
result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output,
 sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2150_c3_9606 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2154_c3_f8a1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2161_c3_374e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2163_c3_f5e2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2158_c7_f092_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2146_l2166_l2158_DUPLICATE_4d74_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2146_l2158_DUPLICATE_1533_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_f480_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2146_l2153_l2158_DUPLICATE_f6f7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_5e95_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2166_l2153_l2158_DUPLICATE_b1a7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5c64_uxn_opcodes_h_l2173_l2142_DUPLICATE_0c4c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2161_c3_374e := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2161_c3_374e;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2163_c3_f5e2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2163_c3_f5e2;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2154_c3_f8a1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2154_c3_f8a1;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2150_c3_9606 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2150_c3_9606;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2153_c11_adc8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2166_c11_c6d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2166_l2153_l2158_DUPLICATE_b1a7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2166_l2153_l2158_DUPLICATE_b1a7_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2146_l2166_l2158_DUPLICATE_4d74 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2146_l2166_l2158_DUPLICATE_4d74_return_output := result.is_sp_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2158_c7_f092_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2146_l2153_l2158_DUPLICATE_f6f7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2146_l2153_l2158_DUPLICATE_f6f7_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_f480 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_f480_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2156_c30_9b72] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_ins;
     sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_x;
     sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output := sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2146_c6_de3d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2158_c11_2195] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_left;
     BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output := BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_5e95 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_5e95_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2146_l2158_DUPLICATE_1533 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2146_l2158_DUPLICATE_1533_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2146_c6_de3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2153_c11_adc8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2158_c11_2195_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2166_c11_c6d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2146_l2158_DUPLICATE_1533_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2146_l2158_DUPLICATE_1533_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2166_l2153_l2158_DUPLICATE_b1a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2166_l2153_l2158_DUPLICATE_b1a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2166_l2153_l2158_DUPLICATE_b1a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2146_l2166_l2158_DUPLICATE_4d74_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2146_l2166_l2158_DUPLICATE_4d74_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2146_l2166_l2158_DUPLICATE_4d74_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_f480_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_f480_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_f480_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_5e95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_5e95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2146_l2166_l2153_DUPLICATE_5e95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2146_l2153_l2158_DUPLICATE_f6f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2146_l2153_l2158_DUPLICATE_f6f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2146_l2153_l2158_DUPLICATE_f6f7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2156_c30_9b72_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2166_c7_a66e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- t8_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     t8_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     t8_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2166_c7_a66e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2166_c7_a66e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2166_c7_a66e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2166_c7_a66e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     -- t8_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2158_c7_f092] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2158_c7_f092_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2153_c7_55d2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2153_c7_55d2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2146_c2_ee74] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output;

     -- Submodule level 5
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5c64_uxn_opcodes_h_l2173_l2142_DUPLICATE_0c4c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5c64_uxn_opcodes_h_l2173_l2142_DUPLICATE_0c4c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5c64(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2146_c2_ee74_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5c64_uxn_opcodes_h_l2173_l2142_DUPLICATE_0c4c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5c64_uxn_opcodes_h_l2173_l2142_DUPLICATE_0c4c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
