-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_929b]
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1162_c2_f867]
signal n8_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_f867]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1162_c2_f867]
signal t8_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1175_c11_dcf7]
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal n8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1175_c7_50c9]
signal t8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1178_c11_6a43]
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal n8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1178_c7_4a57]
signal t8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1181_c11_941b]
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1181_c7_bcac]
signal n8_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1181_c7_bcac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1181_c7_bcac]
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1181_c7_bcac]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1181_c7_bcac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1181_c7_bcac]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1183_c30_0efa]
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1186_c21_52be]
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1186_c21_fdd8]
signal MUX_uxn_opcodes_h_l1186_c21_fdd8_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_fdd8_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_fdd8_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_left,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_right,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output);

-- n8_MUX_uxn_opcodes_h_l1162_c2_f867
n8_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
n8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
n8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- t8_MUX_uxn_opcodes_h_l1162_c2_f867
t8_MUX_uxn_opcodes_h_l1162_c2_f867 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1162_c2_f867_cond,
t8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue,
t8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse,
t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_left,
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_right,
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output);

-- n8_MUX_uxn_opcodes_h_l1175_c7_50c9
n8_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- t8_MUX_uxn_opcodes_h_l1175_c7_50c9
t8_MUX_uxn_opcodes_h_l1175_c7_50c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond,
t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue,
t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse,
t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_left,
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_right,
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output);

-- n8_MUX_uxn_opcodes_h_l1178_c7_4a57
n8_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- t8_MUX_uxn_opcodes_h_l1178_c7_4a57
t8_MUX_uxn_opcodes_h_l1178_c7_4a57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond,
t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue,
t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse,
t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_left,
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_right,
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output);

-- n8_MUX_uxn_opcodes_h_l1181_c7_bcac
n8_MUX_uxn_opcodes_h_l1181_c7_bcac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1181_c7_bcac_cond,
n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue,
n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse,
n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_cond,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa
sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_ins,
sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_x,
sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_y,
sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_left,
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_right,
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output);

-- MUX_uxn_opcodes_h_l1186_c21_fdd8
MUX_uxn_opcodes_h_l1186_c21_fdd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1186_c21_fdd8_cond,
MUX_uxn_opcodes_h_l1186_c21_fdd8_iftrue,
MUX_uxn_opcodes_h_l1186_c21_fdd8_iffalse,
MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output,
 n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output,
 n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output,
 n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output,
 n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output,
 sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output,
 MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_fd67 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_2c04 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_d624 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_9925 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_99ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_467f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_28fd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_2363_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1158_l1190_DUPLICATE_d818_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_2c04 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_2c04;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_d624 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_d624;
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_right := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_right := to_unsigned(3, 2);
     VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_9925 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_9925;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_fd67 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_fd67;
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_929b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_f867_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1183_c30_0efa] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_ins;
     sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_x;
     sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output := sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1186_c21_52be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_left;
     BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output := BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1181_c11_941b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_99ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_99ba_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1178_c11_6a43] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_left;
     BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output := BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_f867_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_f867_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_467f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_467f_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_2363 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_2363_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_28fd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_28fd_return_output := result.is_opc_done;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_f867_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1175_c11_dcf7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_929b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_dcf7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6a43_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_941b_return_output;
     VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_52be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_467f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_467f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_467f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_28fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_28fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_28fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_99ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_99ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1178_l1181_DUPLICATE_99ba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_2363_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_2363_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1178_l1162_l1181_DUPLICATE_88ae_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_f867_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_f867_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_f867_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_f867_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_0efa_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- MUX[uxn_opcodes_h_l1186_c21_fdd8] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1186_c21_fdd8_cond <= VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_cond;
     MUX_uxn_opcodes_h_l1186_c21_fdd8_iftrue <= VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_iftrue;
     MUX_uxn_opcodes_h_l1186_c21_fdd8_iffalse <= VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output := MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- n8_MUX[uxn_opcodes_h_l1181_c7_bcac] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1181_c7_bcac_cond <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_cond;
     n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue;
     n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output := n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1181_c7_bcac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1181_c7_bcac] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1181_c7_bcac] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;

     -- t8_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1181_c7_bcac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue := VAR_MUX_uxn_opcodes_h_l1186_c21_fdd8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1181_c7_bcac] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output := result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;

     -- t8_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- n8_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bcac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     t8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     t8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1178_c7_4a57] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output := result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_4a57_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1175_c7_50c9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- n8_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     n8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     n8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_50c9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_f867] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output := result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1158_l1190_DUPLICATE_d818 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1158_l1190_DUPLICATE_d818_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_f867_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_f867_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1158_l1190_DUPLICATE_d818_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1158_l1190_DUPLICATE_d818_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
