-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity jsr2_0CLK_609876da is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr2_0CLK_609876da;
architecture arch of jsr2_0CLK_609876da is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l773_c6_08cb]
signal BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l773_c2_41c0]
signal t16_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l773_c2_41c0]
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l786_c11_4543]
signal BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l786_c7_c97a]
signal t16_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l786_c7_c97a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l789_c11_eb83]
signal BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l789_c7_3855]
signal t16_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l789_c7_3855]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l791_c3_8319]
signal CONST_SL_8_uxn_opcodes_h_l791_c3_8319_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l792_c30_904a]
signal sp_relative_shift_uxn_opcodes_h_l792_c30_904a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l792_c30_904a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l792_c30_904a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l794_c11_dcc2]
signal BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal t16_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l794_c7_5ea8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l795_c3_9304]
signal BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l802_c11_0a46]
signal BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l802_c7_edcb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l802_c7_edcb]
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l802_c7_edcb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l802_c7_edcb]
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l802_c7_edcb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l802_c7_edcb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l805_c31_cd38]
signal CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output : unsigned(15 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_d736( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.u16_value := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_vram_write := ref_toks_9;
      base.u8_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb
BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_left,
BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_right,
BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output);

-- t16_MUX_uxn_opcodes_h_l773_c2_41c0
t16_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
t16_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
t16_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0
result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0
result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond,
result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543
BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_left,
BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_right,
BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output);

-- t16_MUX_uxn_opcodes_h_l786_c7_c97a
t16_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
t16_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
t16_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a
result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a
result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83
BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_left,
BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_right,
BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output);

-- t16_MUX_uxn_opcodes_h_l789_c7_3855
t16_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l789_c7_3855_cond,
t16_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
t16_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855
result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855
result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output);

-- CONST_SL_8_uxn_opcodes_h_l791_c3_8319
CONST_SL_8_uxn_opcodes_h_l791_c3_8319 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l791_c3_8319_x,
CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output);

-- sp_relative_shift_uxn_opcodes_h_l792_c30_904a
sp_relative_shift_uxn_opcodes_h_l792_c30_904a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l792_c30_904a_ins,
sp_relative_shift_uxn_opcodes_h_l792_c30_904a_x,
sp_relative_shift_uxn_opcodes_h_l792_c30_904a_y,
sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2
BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_left,
BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_right,
BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output);

-- t16_MUX_uxn_opcodes_h_l794_c7_5ea8
t16_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8
result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8
result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l795_c3_9304
BIN_OP_OR_uxn_opcodes_h_l795_c3_9304 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_left,
BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_right,
BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46
BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_left,
BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_right,
BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb
result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond,
result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb
result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond,
result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output);

-- CONST_SR_8_uxn_opcodes_h_l805_c31_cd38
CONST_SR_8_uxn_opcodes_h_l805_c31_cd38 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_x,
CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output,
 t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output,
 t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output,
 t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output,
 CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output,
 sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output,
 t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output,
 BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output,
 CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l778_c3_7990 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l783_c3_166c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l787_c3_ebf4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8319_x : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l799_c3_2eeb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l797_c3_859e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l800_c21_4955_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l803_c3_0f5f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_5f08 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l805_c21_0173_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_9224_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_64ed_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l802_l786_DUPLICATE_d25e_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_8509_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l802_l789_DUPLICATE_bc79_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l769_l811_DUPLICATE_92be_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_5f08 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_5f08;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l803_c3_0f5f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l803_c3_0f5f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l787_c3_ebf4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l787_c3_ebf4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l778_c3_7990 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l778_c3_7990;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l799_c3_2eeb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l799_c3_2eeb;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l783_c3_166c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l783_c3_166c;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l797_c3_859e := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l797_c3_859e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_ins := VAR_ins;
     VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := t16;
     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_8509 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_8509_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l802_l789_DUPLICATE_bc79 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l802_l789_DUPLICATE_bc79_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l773_c6_08cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_9224 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_9224_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l789_c11_eb83] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_left;
     BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output := BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l794_c11_dcc2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_left;
     BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output := BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l805_c31_cd38] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_x <= VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output := CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_64ed LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_64ed_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l773_c2_41c0_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l773_c2_41c0_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l802_l786_DUPLICATE_d25e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l802_l786_DUPLICATE_d25e_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l786_c11_4543] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_left;
     BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output := BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l792_c30_904a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l792_c30_904a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_ins;
     sp_relative_shift_uxn_opcodes_h_l792_c30_904a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_x;
     sp_relative_shift_uxn_opcodes_h_l792_c30_904a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output := sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l800_c21_4955] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l800_c21_4955_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l802_c11_0a46] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_left;
     BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output := BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_08cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_4543_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_eb83_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_dcc2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_0a46_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_8509_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8319_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_8509_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l800_c21_4955_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l802_l786_DUPLICATE_d25e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l802_l786_DUPLICATE_d25e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l802_l794_l789_l786_l773_DUPLICATE_639b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_bd9c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l802_l789_l794_l786_DUPLICATE_477a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_9224_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_9224_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_9224_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_64ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_64ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l789_l794_l786_DUPLICATE_64ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l802_l789_DUPLICATE_bc79_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l802_l789_DUPLICATE_bc79_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l802_l789_l773_l786_DUPLICATE_adb8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l773_c2_41c0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l773_c2_41c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_904a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l802_c7_edcb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l795_c3_9304] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_left;
     BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output := BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l802_c7_edcb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output := result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l802_c7_edcb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l802_c7_edcb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l802_c7_edcb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l805_c21_0173] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l805_c21_0173_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_cd38_return_output);

     -- result_is_vram_write_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l791_c3_8319] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l791_c3_8319_x <= VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8319_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output := CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_9304_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l805_c21_0173_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8319_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- t16_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l802_c7_edcb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output := result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_edcb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_t16_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l794_c7_5ea8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output := result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- t16_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     t16_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     t16_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output := t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_5ea8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- t16_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     t16_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     t16_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l789_c7_3855] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_cond;
     result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output := result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_3855_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_t16_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l786_c7_c97a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output := result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;

     -- t16_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     t16_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     t16_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_c97a_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l773_c2_41c0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output := result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l769_l811_DUPLICATE_92be LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l769_l811_DUPLICATE_92be_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d736(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_41c0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_41c0_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l769_l811_DUPLICATE_92be_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l769_l811_DUPLICATE_92be_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
