-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 134
entity uint8_mux128_0CLK_9347d63d is
port(
 sel : in unsigned(6 downto 0);
 in0 : in unsigned(7 downto 0);
 in1 : in unsigned(7 downto 0);
 in2 : in unsigned(7 downto 0);
 in3 : in unsigned(7 downto 0);
 in4 : in unsigned(7 downto 0);
 in5 : in unsigned(7 downto 0);
 in6 : in unsigned(7 downto 0);
 in7 : in unsigned(7 downto 0);
 in8 : in unsigned(7 downto 0);
 in9 : in unsigned(7 downto 0);
 in10 : in unsigned(7 downto 0);
 in11 : in unsigned(7 downto 0);
 in12 : in unsigned(7 downto 0);
 in13 : in unsigned(7 downto 0);
 in14 : in unsigned(7 downto 0);
 in15 : in unsigned(7 downto 0);
 in16 : in unsigned(7 downto 0);
 in17 : in unsigned(7 downto 0);
 in18 : in unsigned(7 downto 0);
 in19 : in unsigned(7 downto 0);
 in20 : in unsigned(7 downto 0);
 in21 : in unsigned(7 downto 0);
 in22 : in unsigned(7 downto 0);
 in23 : in unsigned(7 downto 0);
 in24 : in unsigned(7 downto 0);
 in25 : in unsigned(7 downto 0);
 in26 : in unsigned(7 downto 0);
 in27 : in unsigned(7 downto 0);
 in28 : in unsigned(7 downto 0);
 in29 : in unsigned(7 downto 0);
 in30 : in unsigned(7 downto 0);
 in31 : in unsigned(7 downto 0);
 in32 : in unsigned(7 downto 0);
 in33 : in unsigned(7 downto 0);
 in34 : in unsigned(7 downto 0);
 in35 : in unsigned(7 downto 0);
 in36 : in unsigned(7 downto 0);
 in37 : in unsigned(7 downto 0);
 in38 : in unsigned(7 downto 0);
 in39 : in unsigned(7 downto 0);
 in40 : in unsigned(7 downto 0);
 in41 : in unsigned(7 downto 0);
 in42 : in unsigned(7 downto 0);
 in43 : in unsigned(7 downto 0);
 in44 : in unsigned(7 downto 0);
 in45 : in unsigned(7 downto 0);
 in46 : in unsigned(7 downto 0);
 in47 : in unsigned(7 downto 0);
 in48 : in unsigned(7 downto 0);
 in49 : in unsigned(7 downto 0);
 in50 : in unsigned(7 downto 0);
 in51 : in unsigned(7 downto 0);
 in52 : in unsigned(7 downto 0);
 in53 : in unsigned(7 downto 0);
 in54 : in unsigned(7 downto 0);
 in55 : in unsigned(7 downto 0);
 in56 : in unsigned(7 downto 0);
 in57 : in unsigned(7 downto 0);
 in58 : in unsigned(7 downto 0);
 in59 : in unsigned(7 downto 0);
 in60 : in unsigned(7 downto 0);
 in61 : in unsigned(7 downto 0);
 in62 : in unsigned(7 downto 0);
 in63 : in unsigned(7 downto 0);
 in64 : in unsigned(7 downto 0);
 in65 : in unsigned(7 downto 0);
 in66 : in unsigned(7 downto 0);
 in67 : in unsigned(7 downto 0);
 in68 : in unsigned(7 downto 0);
 in69 : in unsigned(7 downto 0);
 in70 : in unsigned(7 downto 0);
 in71 : in unsigned(7 downto 0);
 in72 : in unsigned(7 downto 0);
 in73 : in unsigned(7 downto 0);
 in74 : in unsigned(7 downto 0);
 in75 : in unsigned(7 downto 0);
 in76 : in unsigned(7 downto 0);
 in77 : in unsigned(7 downto 0);
 in78 : in unsigned(7 downto 0);
 in79 : in unsigned(7 downto 0);
 in80 : in unsigned(7 downto 0);
 in81 : in unsigned(7 downto 0);
 in82 : in unsigned(7 downto 0);
 in83 : in unsigned(7 downto 0);
 in84 : in unsigned(7 downto 0);
 in85 : in unsigned(7 downto 0);
 in86 : in unsigned(7 downto 0);
 in87 : in unsigned(7 downto 0);
 in88 : in unsigned(7 downto 0);
 in89 : in unsigned(7 downto 0);
 in90 : in unsigned(7 downto 0);
 in91 : in unsigned(7 downto 0);
 in92 : in unsigned(7 downto 0);
 in93 : in unsigned(7 downto 0);
 in94 : in unsigned(7 downto 0);
 in95 : in unsigned(7 downto 0);
 in96 : in unsigned(7 downto 0);
 in97 : in unsigned(7 downto 0);
 in98 : in unsigned(7 downto 0);
 in99 : in unsigned(7 downto 0);
 in100 : in unsigned(7 downto 0);
 in101 : in unsigned(7 downto 0);
 in102 : in unsigned(7 downto 0);
 in103 : in unsigned(7 downto 0);
 in104 : in unsigned(7 downto 0);
 in105 : in unsigned(7 downto 0);
 in106 : in unsigned(7 downto 0);
 in107 : in unsigned(7 downto 0);
 in108 : in unsigned(7 downto 0);
 in109 : in unsigned(7 downto 0);
 in110 : in unsigned(7 downto 0);
 in111 : in unsigned(7 downto 0);
 in112 : in unsigned(7 downto 0);
 in113 : in unsigned(7 downto 0);
 in114 : in unsigned(7 downto 0);
 in115 : in unsigned(7 downto 0);
 in116 : in unsigned(7 downto 0);
 in117 : in unsigned(7 downto 0);
 in118 : in unsigned(7 downto 0);
 in119 : in unsigned(7 downto 0);
 in120 : in unsigned(7 downto 0);
 in121 : in unsigned(7 downto 0);
 in122 : in unsigned(7 downto 0);
 in123 : in unsigned(7 downto 0);
 in124 : in unsigned(7 downto 0);
 in125 : in unsigned(7 downto 0);
 in126 : in unsigned(7 downto 0);
 in127 : in unsigned(7 downto 0);
 return_output : out unsigned(7 downto 0));
end uint8_mux128_0CLK_9347d63d;
architecture arch of uint8_mux128_0CLK_9347d63d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_5094]
signal layer0_node0_MUX_bit_math_h_l18_c3_5094_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_5094_iftrue : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_5094_iffalse : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output : unsigned(7 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_419a]
signal layer0_node1_MUX_bit_math_h_l29_c3_419a_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_419a_iftrue : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_419a_iffalse : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output : unsigned(7 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_195c]
signal layer0_node2_MUX_bit_math_h_l40_c3_195c_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_195c_iftrue : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_195c_iffalse : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output : unsigned(7 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_7a6b]
signal layer0_node3_MUX_bit_math_h_l51_c3_7a6b_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iftrue : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iffalse : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output : unsigned(7 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_1ccf]
signal layer0_node4_MUX_bit_math_h_l62_c3_1ccf_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iftrue : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iffalse : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output : unsigned(7 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_0dd3]
signal layer0_node5_MUX_bit_math_h_l73_c3_0dd3_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iftrue : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iffalse : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output : unsigned(7 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_7e59]
signal layer0_node6_MUX_bit_math_h_l84_c3_7e59_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_7e59_iftrue : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_7e59_iffalse : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output : unsigned(7 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_ffca]
signal layer0_node7_MUX_bit_math_h_l95_c3_ffca_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_ffca_iftrue : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_ffca_iffalse : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output : unsigned(7 downto 0);

-- layer0_node8_MUX[bit_math_h_l106_c3_0c54]
signal layer0_node8_MUX_bit_math_h_l106_c3_0c54_cond : unsigned(0 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_0c54_iftrue : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_0c54_iffalse : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output : unsigned(7 downto 0);

-- layer0_node9_MUX[bit_math_h_l117_c3_521d]
signal layer0_node9_MUX_bit_math_h_l117_c3_521d_cond : unsigned(0 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_521d_iftrue : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_521d_iffalse : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output : unsigned(7 downto 0);

-- layer0_node10_MUX[bit_math_h_l128_c3_74ca]
signal layer0_node10_MUX_bit_math_h_l128_c3_74ca_cond : unsigned(0 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_74ca_iftrue : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_74ca_iffalse : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output : unsigned(7 downto 0);

-- layer0_node11_MUX[bit_math_h_l139_c3_31b7]
signal layer0_node11_MUX_bit_math_h_l139_c3_31b7_cond : unsigned(0 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_31b7_iftrue : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_31b7_iffalse : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output : unsigned(7 downto 0);

-- layer0_node12_MUX[bit_math_h_l150_c3_ce47]
signal layer0_node12_MUX_bit_math_h_l150_c3_ce47_cond : unsigned(0 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_ce47_iftrue : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_ce47_iffalse : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output : unsigned(7 downto 0);

-- layer0_node13_MUX[bit_math_h_l161_c3_76bd]
signal layer0_node13_MUX_bit_math_h_l161_c3_76bd_cond : unsigned(0 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_76bd_iftrue : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_76bd_iffalse : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output : unsigned(7 downto 0);

-- layer0_node14_MUX[bit_math_h_l172_c3_7b21]
signal layer0_node14_MUX_bit_math_h_l172_c3_7b21_cond : unsigned(0 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_7b21_iftrue : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_7b21_iffalse : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output : unsigned(7 downto 0);

-- layer0_node15_MUX[bit_math_h_l183_c3_d015]
signal layer0_node15_MUX_bit_math_h_l183_c3_d015_cond : unsigned(0 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_d015_iftrue : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_d015_iffalse : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output : unsigned(7 downto 0);

-- layer0_node16_MUX[bit_math_h_l194_c3_2677]
signal layer0_node16_MUX_bit_math_h_l194_c3_2677_cond : unsigned(0 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_2677_iftrue : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_2677_iffalse : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output : unsigned(7 downto 0);

-- layer0_node17_MUX[bit_math_h_l205_c3_983c]
signal layer0_node17_MUX_bit_math_h_l205_c3_983c_cond : unsigned(0 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_983c_iftrue : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_983c_iffalse : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output : unsigned(7 downto 0);

-- layer0_node18_MUX[bit_math_h_l216_c3_6aca]
signal layer0_node18_MUX_bit_math_h_l216_c3_6aca_cond : unsigned(0 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_6aca_iftrue : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_6aca_iffalse : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output : unsigned(7 downto 0);

-- layer0_node19_MUX[bit_math_h_l227_c3_1ba6]
signal layer0_node19_MUX_bit_math_h_l227_c3_1ba6_cond : unsigned(0 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iftrue : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iffalse : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output : unsigned(7 downto 0);

-- layer0_node20_MUX[bit_math_h_l238_c3_27b2]
signal layer0_node20_MUX_bit_math_h_l238_c3_27b2_cond : unsigned(0 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_27b2_iftrue : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_27b2_iffalse : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output : unsigned(7 downto 0);

-- layer0_node21_MUX[bit_math_h_l249_c3_c899]
signal layer0_node21_MUX_bit_math_h_l249_c3_c899_cond : unsigned(0 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_c899_iftrue : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_c899_iffalse : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output : unsigned(7 downto 0);

-- layer0_node22_MUX[bit_math_h_l260_c3_0382]
signal layer0_node22_MUX_bit_math_h_l260_c3_0382_cond : unsigned(0 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_0382_iftrue : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_0382_iffalse : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output : unsigned(7 downto 0);

-- layer0_node23_MUX[bit_math_h_l271_c3_93d7]
signal layer0_node23_MUX_bit_math_h_l271_c3_93d7_cond : unsigned(0 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_93d7_iftrue : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_93d7_iffalse : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output : unsigned(7 downto 0);

-- layer0_node24_MUX[bit_math_h_l282_c3_de03]
signal layer0_node24_MUX_bit_math_h_l282_c3_de03_cond : unsigned(0 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_de03_iftrue : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_de03_iffalse : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output : unsigned(7 downto 0);

-- layer0_node25_MUX[bit_math_h_l293_c3_32f2]
signal layer0_node25_MUX_bit_math_h_l293_c3_32f2_cond : unsigned(0 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_32f2_iftrue : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_32f2_iffalse : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output : unsigned(7 downto 0);

-- layer0_node26_MUX[bit_math_h_l304_c3_53c3]
signal layer0_node26_MUX_bit_math_h_l304_c3_53c3_cond : unsigned(0 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_53c3_iftrue : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_53c3_iffalse : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output : unsigned(7 downto 0);

-- layer0_node27_MUX[bit_math_h_l315_c3_e4a1]
signal layer0_node27_MUX_bit_math_h_l315_c3_e4a1_cond : unsigned(0 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iftrue : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iffalse : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output : unsigned(7 downto 0);

-- layer0_node28_MUX[bit_math_h_l326_c3_a3f6]
signal layer0_node28_MUX_bit_math_h_l326_c3_a3f6_cond : unsigned(0 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iftrue : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iffalse : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output : unsigned(7 downto 0);

-- layer0_node29_MUX[bit_math_h_l337_c3_76ce]
signal layer0_node29_MUX_bit_math_h_l337_c3_76ce_cond : unsigned(0 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_76ce_iftrue : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_76ce_iffalse : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output : unsigned(7 downto 0);

-- layer0_node30_MUX[bit_math_h_l348_c3_c538]
signal layer0_node30_MUX_bit_math_h_l348_c3_c538_cond : unsigned(0 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_c538_iftrue : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_c538_iffalse : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output : unsigned(7 downto 0);

-- layer0_node31_MUX[bit_math_h_l359_c3_a259]
signal layer0_node31_MUX_bit_math_h_l359_c3_a259_cond : unsigned(0 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_a259_iftrue : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_a259_iffalse : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output : unsigned(7 downto 0);

-- layer0_node32_MUX[bit_math_h_l370_c3_2900]
signal layer0_node32_MUX_bit_math_h_l370_c3_2900_cond : unsigned(0 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_2900_iftrue : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_2900_iffalse : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output : unsigned(7 downto 0);

-- layer0_node33_MUX[bit_math_h_l381_c3_53ee]
signal layer0_node33_MUX_bit_math_h_l381_c3_53ee_cond : unsigned(0 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_53ee_iftrue : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_53ee_iffalse : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output : unsigned(7 downto 0);

-- layer0_node34_MUX[bit_math_h_l392_c3_e101]
signal layer0_node34_MUX_bit_math_h_l392_c3_e101_cond : unsigned(0 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_e101_iftrue : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_e101_iffalse : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output : unsigned(7 downto 0);

-- layer0_node35_MUX[bit_math_h_l403_c3_00e8]
signal layer0_node35_MUX_bit_math_h_l403_c3_00e8_cond : unsigned(0 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_00e8_iftrue : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_00e8_iffalse : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output : unsigned(7 downto 0);

-- layer0_node36_MUX[bit_math_h_l414_c3_d477]
signal layer0_node36_MUX_bit_math_h_l414_c3_d477_cond : unsigned(0 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_d477_iftrue : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_d477_iffalse : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output : unsigned(7 downto 0);

-- layer0_node37_MUX[bit_math_h_l425_c3_bb07]
signal layer0_node37_MUX_bit_math_h_l425_c3_bb07_cond : unsigned(0 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_bb07_iftrue : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_bb07_iffalse : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output : unsigned(7 downto 0);

-- layer0_node38_MUX[bit_math_h_l436_c3_0345]
signal layer0_node38_MUX_bit_math_h_l436_c3_0345_cond : unsigned(0 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_0345_iftrue : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_0345_iffalse : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output : unsigned(7 downto 0);

-- layer0_node39_MUX[bit_math_h_l447_c3_50eb]
signal layer0_node39_MUX_bit_math_h_l447_c3_50eb_cond : unsigned(0 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_50eb_iftrue : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_50eb_iffalse : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output : unsigned(7 downto 0);

-- layer0_node40_MUX[bit_math_h_l458_c3_0262]
signal layer0_node40_MUX_bit_math_h_l458_c3_0262_cond : unsigned(0 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_0262_iftrue : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_0262_iffalse : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output : unsigned(7 downto 0);

-- layer0_node41_MUX[bit_math_h_l469_c3_4656]
signal layer0_node41_MUX_bit_math_h_l469_c3_4656_cond : unsigned(0 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_4656_iftrue : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_4656_iffalse : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output : unsigned(7 downto 0);

-- layer0_node42_MUX[bit_math_h_l480_c3_45fb]
signal layer0_node42_MUX_bit_math_h_l480_c3_45fb_cond : unsigned(0 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_45fb_iftrue : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_45fb_iffalse : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output : unsigned(7 downto 0);

-- layer0_node43_MUX[bit_math_h_l491_c3_0137]
signal layer0_node43_MUX_bit_math_h_l491_c3_0137_cond : unsigned(0 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_0137_iftrue : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_0137_iffalse : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output : unsigned(7 downto 0);

-- layer0_node44_MUX[bit_math_h_l502_c3_983c]
signal layer0_node44_MUX_bit_math_h_l502_c3_983c_cond : unsigned(0 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_983c_iftrue : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_983c_iffalse : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output : unsigned(7 downto 0);

-- layer0_node45_MUX[bit_math_h_l513_c3_405f]
signal layer0_node45_MUX_bit_math_h_l513_c3_405f_cond : unsigned(0 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_405f_iftrue : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_405f_iffalse : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output : unsigned(7 downto 0);

-- layer0_node46_MUX[bit_math_h_l524_c3_1b28]
signal layer0_node46_MUX_bit_math_h_l524_c3_1b28_cond : unsigned(0 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_1b28_iftrue : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_1b28_iffalse : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output : unsigned(7 downto 0);

-- layer0_node47_MUX[bit_math_h_l535_c3_8ede]
signal layer0_node47_MUX_bit_math_h_l535_c3_8ede_cond : unsigned(0 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_8ede_iftrue : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_8ede_iffalse : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output : unsigned(7 downto 0);

-- layer0_node48_MUX[bit_math_h_l546_c3_f942]
signal layer0_node48_MUX_bit_math_h_l546_c3_f942_cond : unsigned(0 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_f942_iftrue : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_f942_iffalse : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output : unsigned(7 downto 0);

-- layer0_node49_MUX[bit_math_h_l557_c3_44e2]
signal layer0_node49_MUX_bit_math_h_l557_c3_44e2_cond : unsigned(0 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_44e2_iftrue : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_44e2_iffalse : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output : unsigned(7 downto 0);

-- layer0_node50_MUX[bit_math_h_l568_c3_1207]
signal layer0_node50_MUX_bit_math_h_l568_c3_1207_cond : unsigned(0 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_1207_iftrue : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_1207_iffalse : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output : unsigned(7 downto 0);

-- layer0_node51_MUX[bit_math_h_l579_c3_a08f]
signal layer0_node51_MUX_bit_math_h_l579_c3_a08f_cond : unsigned(0 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_a08f_iftrue : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_a08f_iffalse : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output : unsigned(7 downto 0);

-- layer0_node52_MUX[bit_math_h_l590_c3_f2e8]
signal layer0_node52_MUX_bit_math_h_l590_c3_f2e8_cond : unsigned(0 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iftrue : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iffalse : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output : unsigned(7 downto 0);

-- layer0_node53_MUX[bit_math_h_l601_c3_33d0]
signal layer0_node53_MUX_bit_math_h_l601_c3_33d0_cond : unsigned(0 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_33d0_iftrue : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_33d0_iffalse : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output : unsigned(7 downto 0);

-- layer0_node54_MUX[bit_math_h_l612_c3_b44b]
signal layer0_node54_MUX_bit_math_h_l612_c3_b44b_cond : unsigned(0 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_b44b_iftrue : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_b44b_iffalse : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output : unsigned(7 downto 0);

-- layer0_node55_MUX[bit_math_h_l623_c3_0aaf]
signal layer0_node55_MUX_bit_math_h_l623_c3_0aaf_cond : unsigned(0 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iftrue : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iffalse : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output : unsigned(7 downto 0);

-- layer0_node56_MUX[bit_math_h_l634_c3_6313]
signal layer0_node56_MUX_bit_math_h_l634_c3_6313_cond : unsigned(0 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_6313_iftrue : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_6313_iffalse : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output : unsigned(7 downto 0);

-- layer0_node57_MUX[bit_math_h_l645_c3_d8b1]
signal layer0_node57_MUX_bit_math_h_l645_c3_d8b1_cond : unsigned(0 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iftrue : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iffalse : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output : unsigned(7 downto 0);

-- layer0_node58_MUX[bit_math_h_l656_c3_485d]
signal layer0_node58_MUX_bit_math_h_l656_c3_485d_cond : unsigned(0 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_485d_iftrue : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_485d_iffalse : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output : unsigned(7 downto 0);

-- layer0_node59_MUX[bit_math_h_l667_c3_6892]
signal layer0_node59_MUX_bit_math_h_l667_c3_6892_cond : unsigned(0 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_6892_iftrue : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_6892_iffalse : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output : unsigned(7 downto 0);

-- layer0_node60_MUX[bit_math_h_l678_c3_51ce]
signal layer0_node60_MUX_bit_math_h_l678_c3_51ce_cond : unsigned(0 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_51ce_iftrue : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_51ce_iffalse : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output : unsigned(7 downto 0);

-- layer0_node61_MUX[bit_math_h_l689_c3_8d98]
signal layer0_node61_MUX_bit_math_h_l689_c3_8d98_cond : unsigned(0 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_8d98_iftrue : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_8d98_iffalse : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output : unsigned(7 downto 0);

-- layer0_node62_MUX[bit_math_h_l700_c3_9327]
signal layer0_node62_MUX_bit_math_h_l700_c3_9327_cond : unsigned(0 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_9327_iftrue : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_9327_iffalse : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output : unsigned(7 downto 0);

-- layer0_node63_MUX[bit_math_h_l711_c3_c233]
signal layer0_node63_MUX_bit_math_h_l711_c3_c233_cond : unsigned(0 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_c233_iftrue : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_c233_iffalse : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output : unsigned(7 downto 0);

-- layer1_node0_MUX[bit_math_h_l728_c3_cd45]
signal layer1_node0_MUX_bit_math_h_l728_c3_cd45_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_cd45_iftrue : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_cd45_iffalse : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output : unsigned(7 downto 0);

-- layer1_node1_MUX[bit_math_h_l739_c3_e269]
signal layer1_node1_MUX_bit_math_h_l739_c3_e269_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_e269_iftrue : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_e269_iffalse : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output : unsigned(7 downto 0);

-- layer1_node2_MUX[bit_math_h_l750_c3_5aa6]
signal layer1_node2_MUX_bit_math_h_l750_c3_5aa6_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iftrue : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iffalse : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output : unsigned(7 downto 0);

-- layer1_node3_MUX[bit_math_h_l761_c3_850a]
signal layer1_node3_MUX_bit_math_h_l761_c3_850a_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_850a_iftrue : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_850a_iffalse : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output : unsigned(7 downto 0);

-- layer1_node4_MUX[bit_math_h_l772_c3_a071]
signal layer1_node4_MUX_bit_math_h_l772_c3_a071_cond : unsigned(0 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_a071_iftrue : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_a071_iffalse : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output : unsigned(7 downto 0);

-- layer1_node5_MUX[bit_math_h_l783_c3_9883]
signal layer1_node5_MUX_bit_math_h_l783_c3_9883_cond : unsigned(0 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_9883_iftrue : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_9883_iffalse : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output : unsigned(7 downto 0);

-- layer1_node6_MUX[bit_math_h_l794_c3_cf43]
signal layer1_node6_MUX_bit_math_h_l794_c3_cf43_cond : unsigned(0 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_cf43_iftrue : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_cf43_iffalse : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output : unsigned(7 downto 0);

-- layer1_node7_MUX[bit_math_h_l805_c3_c99c]
signal layer1_node7_MUX_bit_math_h_l805_c3_c99c_cond : unsigned(0 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_c99c_iftrue : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_c99c_iffalse : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output : unsigned(7 downto 0);

-- layer1_node8_MUX[bit_math_h_l816_c3_fa37]
signal layer1_node8_MUX_bit_math_h_l816_c3_fa37_cond : unsigned(0 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_fa37_iftrue : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_fa37_iffalse : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output : unsigned(7 downto 0);

-- layer1_node9_MUX[bit_math_h_l827_c3_d6c2]
signal layer1_node9_MUX_bit_math_h_l827_c3_d6c2_cond : unsigned(0 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iftrue : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iffalse : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output : unsigned(7 downto 0);

-- layer1_node10_MUX[bit_math_h_l838_c3_7eb8]
signal layer1_node10_MUX_bit_math_h_l838_c3_7eb8_cond : unsigned(0 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iftrue : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iffalse : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output : unsigned(7 downto 0);

-- layer1_node11_MUX[bit_math_h_l849_c3_2cb0]
signal layer1_node11_MUX_bit_math_h_l849_c3_2cb0_cond : unsigned(0 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iftrue : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iffalse : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output : unsigned(7 downto 0);

-- layer1_node12_MUX[bit_math_h_l860_c3_32ef]
signal layer1_node12_MUX_bit_math_h_l860_c3_32ef_cond : unsigned(0 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_32ef_iftrue : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_32ef_iffalse : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output : unsigned(7 downto 0);

-- layer1_node13_MUX[bit_math_h_l871_c3_c37d]
signal layer1_node13_MUX_bit_math_h_l871_c3_c37d_cond : unsigned(0 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_c37d_iftrue : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_c37d_iffalse : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output : unsigned(7 downto 0);

-- layer1_node14_MUX[bit_math_h_l882_c3_3e12]
signal layer1_node14_MUX_bit_math_h_l882_c3_3e12_cond : unsigned(0 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_3e12_iftrue : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_3e12_iffalse : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output : unsigned(7 downto 0);

-- layer1_node15_MUX[bit_math_h_l893_c3_5e2b]
signal layer1_node15_MUX_bit_math_h_l893_c3_5e2b_cond : unsigned(0 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iftrue : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iffalse : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output : unsigned(7 downto 0);

-- layer1_node16_MUX[bit_math_h_l904_c3_234e]
signal layer1_node16_MUX_bit_math_h_l904_c3_234e_cond : unsigned(0 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_234e_iftrue : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_234e_iffalse : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output : unsigned(7 downto 0);

-- layer1_node17_MUX[bit_math_h_l915_c3_90a2]
signal layer1_node17_MUX_bit_math_h_l915_c3_90a2_cond : unsigned(0 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_90a2_iftrue : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_90a2_iffalse : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output : unsigned(7 downto 0);

-- layer1_node18_MUX[bit_math_h_l926_c3_ecc8]
signal layer1_node18_MUX_bit_math_h_l926_c3_ecc8_cond : unsigned(0 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iftrue : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iffalse : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output : unsigned(7 downto 0);

-- layer1_node19_MUX[bit_math_h_l937_c3_7211]
signal layer1_node19_MUX_bit_math_h_l937_c3_7211_cond : unsigned(0 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_7211_iftrue : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_7211_iffalse : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output : unsigned(7 downto 0);

-- layer1_node20_MUX[bit_math_h_l948_c3_2d00]
signal layer1_node20_MUX_bit_math_h_l948_c3_2d00_cond : unsigned(0 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2d00_iftrue : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2d00_iffalse : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output : unsigned(7 downto 0);

-- layer1_node21_MUX[bit_math_h_l959_c3_f682]
signal layer1_node21_MUX_bit_math_h_l959_c3_f682_cond : unsigned(0 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_f682_iftrue : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_f682_iffalse : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output : unsigned(7 downto 0);

-- layer1_node22_MUX[bit_math_h_l970_c3_8998]
signal layer1_node22_MUX_bit_math_h_l970_c3_8998_cond : unsigned(0 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_8998_iftrue : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_8998_iffalse : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output : unsigned(7 downto 0);

-- layer1_node23_MUX[bit_math_h_l981_c3_102a]
signal layer1_node23_MUX_bit_math_h_l981_c3_102a_cond : unsigned(0 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_102a_iftrue : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_102a_iffalse : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output : unsigned(7 downto 0);

-- layer1_node24_MUX[bit_math_h_l992_c3_9fd6]
signal layer1_node24_MUX_bit_math_h_l992_c3_9fd6_cond : unsigned(0 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iftrue : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iffalse : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output : unsigned(7 downto 0);

-- layer1_node25_MUX[bit_math_h_l1003_c3_271e]
signal layer1_node25_MUX_bit_math_h_l1003_c3_271e_cond : unsigned(0 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_271e_iftrue : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_271e_iffalse : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output : unsigned(7 downto 0);

-- layer1_node26_MUX[bit_math_h_l1014_c3_1e7d]
signal layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_cond : unsigned(0 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iftrue : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iffalse : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output : unsigned(7 downto 0);

-- layer1_node27_MUX[bit_math_h_l1025_c3_46dd]
signal layer1_node27_MUX_bit_math_h_l1025_c3_46dd_cond : unsigned(0 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iftrue : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iffalse : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output : unsigned(7 downto 0);

-- layer1_node28_MUX[bit_math_h_l1036_c3_4035]
signal layer1_node28_MUX_bit_math_h_l1036_c3_4035_cond : unsigned(0 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_4035_iftrue : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_4035_iffalse : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output : unsigned(7 downto 0);

-- layer1_node29_MUX[bit_math_h_l1047_c3_3314]
signal layer1_node29_MUX_bit_math_h_l1047_c3_3314_cond : unsigned(0 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_3314_iftrue : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_3314_iffalse : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output : unsigned(7 downto 0);

-- layer1_node30_MUX[bit_math_h_l1058_c3_6a5f]
signal layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_cond : unsigned(0 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iftrue : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iffalse : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output : unsigned(7 downto 0);

-- layer1_node31_MUX[bit_math_h_l1069_c3_5488]
signal layer1_node31_MUX_bit_math_h_l1069_c3_5488_cond : unsigned(0 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_5488_iftrue : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_5488_iffalse : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output : unsigned(7 downto 0);

-- layer2_node0_MUX[bit_math_h_l1086_c3_74df]
signal layer2_node0_MUX_bit_math_h_l1086_c3_74df_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_74df_iftrue : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_74df_iffalse : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output : unsigned(7 downto 0);

-- layer2_node1_MUX[bit_math_h_l1097_c3_4739]
signal layer2_node1_MUX_bit_math_h_l1097_c3_4739_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_4739_iftrue : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_4739_iffalse : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output : unsigned(7 downto 0);

-- layer2_node2_MUX[bit_math_h_l1108_c3_c83e]
signal layer2_node2_MUX_bit_math_h_l1108_c3_c83e_cond : unsigned(0 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iftrue : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iffalse : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output : unsigned(7 downto 0);

-- layer2_node3_MUX[bit_math_h_l1119_c3_1d4a]
signal layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_cond : unsigned(0 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iftrue : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iffalse : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output : unsigned(7 downto 0);

-- layer2_node4_MUX[bit_math_h_l1130_c3_d0b7]
signal layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_cond : unsigned(0 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iftrue : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iffalse : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output : unsigned(7 downto 0);

-- layer2_node5_MUX[bit_math_h_l1141_c3_a33d]
signal layer2_node5_MUX_bit_math_h_l1141_c3_a33d_cond : unsigned(0 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iftrue : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iffalse : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output : unsigned(7 downto 0);

-- layer2_node6_MUX[bit_math_h_l1152_c3_403d]
signal layer2_node6_MUX_bit_math_h_l1152_c3_403d_cond : unsigned(0 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_403d_iftrue : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_403d_iffalse : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output : unsigned(7 downto 0);

-- layer2_node7_MUX[bit_math_h_l1163_c3_f8a3]
signal layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_cond : unsigned(0 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iftrue : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iffalse : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output : unsigned(7 downto 0);

-- layer2_node8_MUX[bit_math_h_l1174_c3_51d4]
signal layer2_node8_MUX_bit_math_h_l1174_c3_51d4_cond : unsigned(0 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iftrue : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iffalse : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output : unsigned(7 downto 0);

-- layer2_node9_MUX[bit_math_h_l1185_c3_30b5]
signal layer2_node9_MUX_bit_math_h_l1185_c3_30b5_cond : unsigned(0 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iftrue : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iffalse : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output : unsigned(7 downto 0);

-- layer2_node10_MUX[bit_math_h_l1196_c3_6142]
signal layer2_node10_MUX_bit_math_h_l1196_c3_6142_cond : unsigned(0 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_6142_iftrue : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_6142_iffalse : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output : unsigned(7 downto 0);

-- layer2_node11_MUX[bit_math_h_l1207_c3_17d4]
signal layer2_node11_MUX_bit_math_h_l1207_c3_17d4_cond : unsigned(0 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iftrue : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iffalse : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output : unsigned(7 downto 0);

-- layer2_node12_MUX[bit_math_h_l1218_c3_74f5]
signal layer2_node12_MUX_bit_math_h_l1218_c3_74f5_cond : unsigned(0 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iftrue : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iffalse : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output : unsigned(7 downto 0);

-- layer2_node13_MUX[bit_math_h_l1229_c3_af85]
signal layer2_node13_MUX_bit_math_h_l1229_c3_af85_cond : unsigned(0 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_af85_iftrue : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_af85_iffalse : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output : unsigned(7 downto 0);

-- layer2_node14_MUX[bit_math_h_l1240_c3_0287]
signal layer2_node14_MUX_bit_math_h_l1240_c3_0287_cond : unsigned(0 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_0287_iftrue : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_0287_iffalse : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output : unsigned(7 downto 0);

-- layer2_node15_MUX[bit_math_h_l1251_c3_a113]
signal layer2_node15_MUX_bit_math_h_l1251_c3_a113_cond : unsigned(0 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_a113_iftrue : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_a113_iffalse : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output : unsigned(7 downto 0);

-- layer3_node0_MUX[bit_math_h_l1268_c3_1d33]
signal layer3_node0_MUX_bit_math_h_l1268_c3_1d33_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iftrue : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iffalse : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output : unsigned(7 downto 0);

-- layer3_node1_MUX[bit_math_h_l1279_c3_ca08]
signal layer3_node1_MUX_bit_math_h_l1279_c3_ca08_cond : unsigned(0 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iftrue : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iffalse : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output : unsigned(7 downto 0);

-- layer3_node2_MUX[bit_math_h_l1290_c3_581b]
signal layer3_node2_MUX_bit_math_h_l1290_c3_581b_cond : unsigned(0 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_581b_iftrue : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_581b_iffalse : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output : unsigned(7 downto 0);

-- layer3_node3_MUX[bit_math_h_l1301_c3_778a]
signal layer3_node3_MUX_bit_math_h_l1301_c3_778a_cond : unsigned(0 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_778a_iftrue : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_778a_iffalse : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output : unsigned(7 downto 0);

-- layer3_node4_MUX[bit_math_h_l1312_c3_9af8]
signal layer3_node4_MUX_bit_math_h_l1312_c3_9af8_cond : unsigned(0 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iftrue : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iffalse : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output : unsigned(7 downto 0);

-- layer3_node5_MUX[bit_math_h_l1323_c3_8487]
signal layer3_node5_MUX_bit_math_h_l1323_c3_8487_cond : unsigned(0 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_8487_iftrue : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_8487_iffalse : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output : unsigned(7 downto 0);

-- layer3_node6_MUX[bit_math_h_l1334_c3_d703]
signal layer3_node6_MUX_bit_math_h_l1334_c3_d703_cond : unsigned(0 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_d703_iftrue : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_d703_iffalse : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output : unsigned(7 downto 0);

-- layer3_node7_MUX[bit_math_h_l1345_c3_ae83]
signal layer3_node7_MUX_bit_math_h_l1345_c3_ae83_cond : unsigned(0 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iftrue : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iffalse : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output : unsigned(7 downto 0);

-- layer4_node0_MUX[bit_math_h_l1362_c3_0390]
signal layer4_node0_MUX_bit_math_h_l1362_c3_0390_cond : unsigned(0 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_0390_iftrue : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_0390_iffalse : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output : unsigned(7 downto 0);

-- layer4_node1_MUX[bit_math_h_l1373_c3_27d5]
signal layer4_node1_MUX_bit_math_h_l1373_c3_27d5_cond : unsigned(0 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iftrue : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iffalse : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output : unsigned(7 downto 0);

-- layer4_node2_MUX[bit_math_h_l1384_c3_2032]
signal layer4_node2_MUX_bit_math_h_l1384_c3_2032_cond : unsigned(0 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_2032_iftrue : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_2032_iffalse : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output : unsigned(7 downto 0);

-- layer4_node3_MUX[bit_math_h_l1395_c3_ef44]
signal layer4_node3_MUX_bit_math_h_l1395_c3_ef44_cond : unsigned(0 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iftrue : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iffalse : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output : unsigned(7 downto 0);

-- layer5_node0_MUX[bit_math_h_l1412_c3_1733]
signal layer5_node0_MUX_bit_math_h_l1412_c3_1733_cond : unsigned(0 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_1733_iftrue : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_1733_iffalse : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output : unsigned(7 downto 0);

-- layer5_node1_MUX[bit_math_h_l1423_c3_54e8]
signal layer5_node1_MUX_bit_math_h_l1423_c3_54e8_cond : unsigned(0 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iftrue : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iffalse : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output : unsigned(7 downto 0);

-- layer6_node0_MUX[bit_math_h_l1440_c3_c11f]
signal layer6_node0_MUX_bit_math_h_l1440_c3_c11f_cond : unsigned(0 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iftrue : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iffalse : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output : unsigned(7 downto 0);

function uint7_0_0( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint7_1_1( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint7_2_2( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint7_3_3( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;

function uint7_4_4( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(4- i);
      end loop;
return return_output;
end function;

function uint7_5_5( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(5- i);
      end loop;
return return_output;
end function;

function uint7_6_6( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(6- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_5094
layer0_node0_MUX_bit_math_h_l18_c3_5094 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_5094_cond,
layer0_node0_MUX_bit_math_h_l18_c3_5094_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_5094_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_419a
layer0_node1_MUX_bit_math_h_l29_c3_419a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_419a_cond,
layer0_node1_MUX_bit_math_h_l29_c3_419a_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_419a_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_195c
layer0_node2_MUX_bit_math_h_l40_c3_195c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_195c_cond,
layer0_node2_MUX_bit_math_h_l40_c3_195c_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_195c_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_7a6b
layer0_node3_MUX_bit_math_h_l51_c3_7a6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_7a6b_cond,
layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_1ccf
layer0_node4_MUX_bit_math_h_l62_c3_1ccf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_1ccf_cond,
layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_0dd3
layer0_node5_MUX_bit_math_h_l73_c3_0dd3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_0dd3_cond,
layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_7e59
layer0_node6_MUX_bit_math_h_l84_c3_7e59 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_7e59_cond,
layer0_node6_MUX_bit_math_h_l84_c3_7e59_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_7e59_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_ffca
layer0_node7_MUX_bit_math_h_l95_c3_ffca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_ffca_cond,
layer0_node7_MUX_bit_math_h_l95_c3_ffca_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_ffca_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output);

-- layer0_node8_MUX_bit_math_h_l106_c3_0c54
layer0_node8_MUX_bit_math_h_l106_c3_0c54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node8_MUX_bit_math_h_l106_c3_0c54_cond,
layer0_node8_MUX_bit_math_h_l106_c3_0c54_iftrue,
layer0_node8_MUX_bit_math_h_l106_c3_0c54_iffalse,
layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output);

-- layer0_node9_MUX_bit_math_h_l117_c3_521d
layer0_node9_MUX_bit_math_h_l117_c3_521d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node9_MUX_bit_math_h_l117_c3_521d_cond,
layer0_node9_MUX_bit_math_h_l117_c3_521d_iftrue,
layer0_node9_MUX_bit_math_h_l117_c3_521d_iffalse,
layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output);

-- layer0_node10_MUX_bit_math_h_l128_c3_74ca
layer0_node10_MUX_bit_math_h_l128_c3_74ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node10_MUX_bit_math_h_l128_c3_74ca_cond,
layer0_node10_MUX_bit_math_h_l128_c3_74ca_iftrue,
layer0_node10_MUX_bit_math_h_l128_c3_74ca_iffalse,
layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output);

-- layer0_node11_MUX_bit_math_h_l139_c3_31b7
layer0_node11_MUX_bit_math_h_l139_c3_31b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node11_MUX_bit_math_h_l139_c3_31b7_cond,
layer0_node11_MUX_bit_math_h_l139_c3_31b7_iftrue,
layer0_node11_MUX_bit_math_h_l139_c3_31b7_iffalse,
layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output);

-- layer0_node12_MUX_bit_math_h_l150_c3_ce47
layer0_node12_MUX_bit_math_h_l150_c3_ce47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node12_MUX_bit_math_h_l150_c3_ce47_cond,
layer0_node12_MUX_bit_math_h_l150_c3_ce47_iftrue,
layer0_node12_MUX_bit_math_h_l150_c3_ce47_iffalse,
layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output);

-- layer0_node13_MUX_bit_math_h_l161_c3_76bd
layer0_node13_MUX_bit_math_h_l161_c3_76bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node13_MUX_bit_math_h_l161_c3_76bd_cond,
layer0_node13_MUX_bit_math_h_l161_c3_76bd_iftrue,
layer0_node13_MUX_bit_math_h_l161_c3_76bd_iffalse,
layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output);

-- layer0_node14_MUX_bit_math_h_l172_c3_7b21
layer0_node14_MUX_bit_math_h_l172_c3_7b21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node14_MUX_bit_math_h_l172_c3_7b21_cond,
layer0_node14_MUX_bit_math_h_l172_c3_7b21_iftrue,
layer0_node14_MUX_bit_math_h_l172_c3_7b21_iffalse,
layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output);

-- layer0_node15_MUX_bit_math_h_l183_c3_d015
layer0_node15_MUX_bit_math_h_l183_c3_d015 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node15_MUX_bit_math_h_l183_c3_d015_cond,
layer0_node15_MUX_bit_math_h_l183_c3_d015_iftrue,
layer0_node15_MUX_bit_math_h_l183_c3_d015_iffalse,
layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output);

-- layer0_node16_MUX_bit_math_h_l194_c3_2677
layer0_node16_MUX_bit_math_h_l194_c3_2677 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node16_MUX_bit_math_h_l194_c3_2677_cond,
layer0_node16_MUX_bit_math_h_l194_c3_2677_iftrue,
layer0_node16_MUX_bit_math_h_l194_c3_2677_iffalse,
layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output);

-- layer0_node17_MUX_bit_math_h_l205_c3_983c
layer0_node17_MUX_bit_math_h_l205_c3_983c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node17_MUX_bit_math_h_l205_c3_983c_cond,
layer0_node17_MUX_bit_math_h_l205_c3_983c_iftrue,
layer0_node17_MUX_bit_math_h_l205_c3_983c_iffalse,
layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output);

-- layer0_node18_MUX_bit_math_h_l216_c3_6aca
layer0_node18_MUX_bit_math_h_l216_c3_6aca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node18_MUX_bit_math_h_l216_c3_6aca_cond,
layer0_node18_MUX_bit_math_h_l216_c3_6aca_iftrue,
layer0_node18_MUX_bit_math_h_l216_c3_6aca_iffalse,
layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output);

-- layer0_node19_MUX_bit_math_h_l227_c3_1ba6
layer0_node19_MUX_bit_math_h_l227_c3_1ba6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node19_MUX_bit_math_h_l227_c3_1ba6_cond,
layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iftrue,
layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iffalse,
layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output);

-- layer0_node20_MUX_bit_math_h_l238_c3_27b2
layer0_node20_MUX_bit_math_h_l238_c3_27b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node20_MUX_bit_math_h_l238_c3_27b2_cond,
layer0_node20_MUX_bit_math_h_l238_c3_27b2_iftrue,
layer0_node20_MUX_bit_math_h_l238_c3_27b2_iffalse,
layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output);

-- layer0_node21_MUX_bit_math_h_l249_c3_c899
layer0_node21_MUX_bit_math_h_l249_c3_c899 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node21_MUX_bit_math_h_l249_c3_c899_cond,
layer0_node21_MUX_bit_math_h_l249_c3_c899_iftrue,
layer0_node21_MUX_bit_math_h_l249_c3_c899_iffalse,
layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output);

-- layer0_node22_MUX_bit_math_h_l260_c3_0382
layer0_node22_MUX_bit_math_h_l260_c3_0382 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node22_MUX_bit_math_h_l260_c3_0382_cond,
layer0_node22_MUX_bit_math_h_l260_c3_0382_iftrue,
layer0_node22_MUX_bit_math_h_l260_c3_0382_iffalse,
layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output);

-- layer0_node23_MUX_bit_math_h_l271_c3_93d7
layer0_node23_MUX_bit_math_h_l271_c3_93d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node23_MUX_bit_math_h_l271_c3_93d7_cond,
layer0_node23_MUX_bit_math_h_l271_c3_93d7_iftrue,
layer0_node23_MUX_bit_math_h_l271_c3_93d7_iffalse,
layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output);

-- layer0_node24_MUX_bit_math_h_l282_c3_de03
layer0_node24_MUX_bit_math_h_l282_c3_de03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node24_MUX_bit_math_h_l282_c3_de03_cond,
layer0_node24_MUX_bit_math_h_l282_c3_de03_iftrue,
layer0_node24_MUX_bit_math_h_l282_c3_de03_iffalse,
layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output);

-- layer0_node25_MUX_bit_math_h_l293_c3_32f2
layer0_node25_MUX_bit_math_h_l293_c3_32f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node25_MUX_bit_math_h_l293_c3_32f2_cond,
layer0_node25_MUX_bit_math_h_l293_c3_32f2_iftrue,
layer0_node25_MUX_bit_math_h_l293_c3_32f2_iffalse,
layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output);

-- layer0_node26_MUX_bit_math_h_l304_c3_53c3
layer0_node26_MUX_bit_math_h_l304_c3_53c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node26_MUX_bit_math_h_l304_c3_53c3_cond,
layer0_node26_MUX_bit_math_h_l304_c3_53c3_iftrue,
layer0_node26_MUX_bit_math_h_l304_c3_53c3_iffalse,
layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output);

-- layer0_node27_MUX_bit_math_h_l315_c3_e4a1
layer0_node27_MUX_bit_math_h_l315_c3_e4a1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node27_MUX_bit_math_h_l315_c3_e4a1_cond,
layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iftrue,
layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iffalse,
layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output);

-- layer0_node28_MUX_bit_math_h_l326_c3_a3f6
layer0_node28_MUX_bit_math_h_l326_c3_a3f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node28_MUX_bit_math_h_l326_c3_a3f6_cond,
layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iftrue,
layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iffalse,
layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output);

-- layer0_node29_MUX_bit_math_h_l337_c3_76ce
layer0_node29_MUX_bit_math_h_l337_c3_76ce : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node29_MUX_bit_math_h_l337_c3_76ce_cond,
layer0_node29_MUX_bit_math_h_l337_c3_76ce_iftrue,
layer0_node29_MUX_bit_math_h_l337_c3_76ce_iffalse,
layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output);

-- layer0_node30_MUX_bit_math_h_l348_c3_c538
layer0_node30_MUX_bit_math_h_l348_c3_c538 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node30_MUX_bit_math_h_l348_c3_c538_cond,
layer0_node30_MUX_bit_math_h_l348_c3_c538_iftrue,
layer0_node30_MUX_bit_math_h_l348_c3_c538_iffalse,
layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output);

-- layer0_node31_MUX_bit_math_h_l359_c3_a259
layer0_node31_MUX_bit_math_h_l359_c3_a259 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node31_MUX_bit_math_h_l359_c3_a259_cond,
layer0_node31_MUX_bit_math_h_l359_c3_a259_iftrue,
layer0_node31_MUX_bit_math_h_l359_c3_a259_iffalse,
layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output);

-- layer0_node32_MUX_bit_math_h_l370_c3_2900
layer0_node32_MUX_bit_math_h_l370_c3_2900 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node32_MUX_bit_math_h_l370_c3_2900_cond,
layer0_node32_MUX_bit_math_h_l370_c3_2900_iftrue,
layer0_node32_MUX_bit_math_h_l370_c3_2900_iffalse,
layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output);

-- layer0_node33_MUX_bit_math_h_l381_c3_53ee
layer0_node33_MUX_bit_math_h_l381_c3_53ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node33_MUX_bit_math_h_l381_c3_53ee_cond,
layer0_node33_MUX_bit_math_h_l381_c3_53ee_iftrue,
layer0_node33_MUX_bit_math_h_l381_c3_53ee_iffalse,
layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output);

-- layer0_node34_MUX_bit_math_h_l392_c3_e101
layer0_node34_MUX_bit_math_h_l392_c3_e101 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node34_MUX_bit_math_h_l392_c3_e101_cond,
layer0_node34_MUX_bit_math_h_l392_c3_e101_iftrue,
layer0_node34_MUX_bit_math_h_l392_c3_e101_iffalse,
layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output);

-- layer0_node35_MUX_bit_math_h_l403_c3_00e8
layer0_node35_MUX_bit_math_h_l403_c3_00e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node35_MUX_bit_math_h_l403_c3_00e8_cond,
layer0_node35_MUX_bit_math_h_l403_c3_00e8_iftrue,
layer0_node35_MUX_bit_math_h_l403_c3_00e8_iffalse,
layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output);

-- layer0_node36_MUX_bit_math_h_l414_c3_d477
layer0_node36_MUX_bit_math_h_l414_c3_d477 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node36_MUX_bit_math_h_l414_c3_d477_cond,
layer0_node36_MUX_bit_math_h_l414_c3_d477_iftrue,
layer0_node36_MUX_bit_math_h_l414_c3_d477_iffalse,
layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output);

-- layer0_node37_MUX_bit_math_h_l425_c3_bb07
layer0_node37_MUX_bit_math_h_l425_c3_bb07 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node37_MUX_bit_math_h_l425_c3_bb07_cond,
layer0_node37_MUX_bit_math_h_l425_c3_bb07_iftrue,
layer0_node37_MUX_bit_math_h_l425_c3_bb07_iffalse,
layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output);

-- layer0_node38_MUX_bit_math_h_l436_c3_0345
layer0_node38_MUX_bit_math_h_l436_c3_0345 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node38_MUX_bit_math_h_l436_c3_0345_cond,
layer0_node38_MUX_bit_math_h_l436_c3_0345_iftrue,
layer0_node38_MUX_bit_math_h_l436_c3_0345_iffalse,
layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output);

-- layer0_node39_MUX_bit_math_h_l447_c3_50eb
layer0_node39_MUX_bit_math_h_l447_c3_50eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node39_MUX_bit_math_h_l447_c3_50eb_cond,
layer0_node39_MUX_bit_math_h_l447_c3_50eb_iftrue,
layer0_node39_MUX_bit_math_h_l447_c3_50eb_iffalse,
layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output);

-- layer0_node40_MUX_bit_math_h_l458_c3_0262
layer0_node40_MUX_bit_math_h_l458_c3_0262 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node40_MUX_bit_math_h_l458_c3_0262_cond,
layer0_node40_MUX_bit_math_h_l458_c3_0262_iftrue,
layer0_node40_MUX_bit_math_h_l458_c3_0262_iffalse,
layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output);

-- layer0_node41_MUX_bit_math_h_l469_c3_4656
layer0_node41_MUX_bit_math_h_l469_c3_4656 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node41_MUX_bit_math_h_l469_c3_4656_cond,
layer0_node41_MUX_bit_math_h_l469_c3_4656_iftrue,
layer0_node41_MUX_bit_math_h_l469_c3_4656_iffalse,
layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output);

-- layer0_node42_MUX_bit_math_h_l480_c3_45fb
layer0_node42_MUX_bit_math_h_l480_c3_45fb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node42_MUX_bit_math_h_l480_c3_45fb_cond,
layer0_node42_MUX_bit_math_h_l480_c3_45fb_iftrue,
layer0_node42_MUX_bit_math_h_l480_c3_45fb_iffalse,
layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output);

-- layer0_node43_MUX_bit_math_h_l491_c3_0137
layer0_node43_MUX_bit_math_h_l491_c3_0137 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node43_MUX_bit_math_h_l491_c3_0137_cond,
layer0_node43_MUX_bit_math_h_l491_c3_0137_iftrue,
layer0_node43_MUX_bit_math_h_l491_c3_0137_iffalse,
layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output);

-- layer0_node44_MUX_bit_math_h_l502_c3_983c
layer0_node44_MUX_bit_math_h_l502_c3_983c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node44_MUX_bit_math_h_l502_c3_983c_cond,
layer0_node44_MUX_bit_math_h_l502_c3_983c_iftrue,
layer0_node44_MUX_bit_math_h_l502_c3_983c_iffalse,
layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output);

-- layer0_node45_MUX_bit_math_h_l513_c3_405f
layer0_node45_MUX_bit_math_h_l513_c3_405f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node45_MUX_bit_math_h_l513_c3_405f_cond,
layer0_node45_MUX_bit_math_h_l513_c3_405f_iftrue,
layer0_node45_MUX_bit_math_h_l513_c3_405f_iffalse,
layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output);

-- layer0_node46_MUX_bit_math_h_l524_c3_1b28
layer0_node46_MUX_bit_math_h_l524_c3_1b28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node46_MUX_bit_math_h_l524_c3_1b28_cond,
layer0_node46_MUX_bit_math_h_l524_c3_1b28_iftrue,
layer0_node46_MUX_bit_math_h_l524_c3_1b28_iffalse,
layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output);

-- layer0_node47_MUX_bit_math_h_l535_c3_8ede
layer0_node47_MUX_bit_math_h_l535_c3_8ede : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node47_MUX_bit_math_h_l535_c3_8ede_cond,
layer0_node47_MUX_bit_math_h_l535_c3_8ede_iftrue,
layer0_node47_MUX_bit_math_h_l535_c3_8ede_iffalse,
layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output);

-- layer0_node48_MUX_bit_math_h_l546_c3_f942
layer0_node48_MUX_bit_math_h_l546_c3_f942 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node48_MUX_bit_math_h_l546_c3_f942_cond,
layer0_node48_MUX_bit_math_h_l546_c3_f942_iftrue,
layer0_node48_MUX_bit_math_h_l546_c3_f942_iffalse,
layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output);

-- layer0_node49_MUX_bit_math_h_l557_c3_44e2
layer0_node49_MUX_bit_math_h_l557_c3_44e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node49_MUX_bit_math_h_l557_c3_44e2_cond,
layer0_node49_MUX_bit_math_h_l557_c3_44e2_iftrue,
layer0_node49_MUX_bit_math_h_l557_c3_44e2_iffalse,
layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output);

-- layer0_node50_MUX_bit_math_h_l568_c3_1207
layer0_node50_MUX_bit_math_h_l568_c3_1207 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node50_MUX_bit_math_h_l568_c3_1207_cond,
layer0_node50_MUX_bit_math_h_l568_c3_1207_iftrue,
layer0_node50_MUX_bit_math_h_l568_c3_1207_iffalse,
layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output);

-- layer0_node51_MUX_bit_math_h_l579_c3_a08f
layer0_node51_MUX_bit_math_h_l579_c3_a08f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node51_MUX_bit_math_h_l579_c3_a08f_cond,
layer0_node51_MUX_bit_math_h_l579_c3_a08f_iftrue,
layer0_node51_MUX_bit_math_h_l579_c3_a08f_iffalse,
layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output);

-- layer0_node52_MUX_bit_math_h_l590_c3_f2e8
layer0_node52_MUX_bit_math_h_l590_c3_f2e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node52_MUX_bit_math_h_l590_c3_f2e8_cond,
layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iftrue,
layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iffalse,
layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output);

-- layer0_node53_MUX_bit_math_h_l601_c3_33d0
layer0_node53_MUX_bit_math_h_l601_c3_33d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node53_MUX_bit_math_h_l601_c3_33d0_cond,
layer0_node53_MUX_bit_math_h_l601_c3_33d0_iftrue,
layer0_node53_MUX_bit_math_h_l601_c3_33d0_iffalse,
layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output);

-- layer0_node54_MUX_bit_math_h_l612_c3_b44b
layer0_node54_MUX_bit_math_h_l612_c3_b44b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node54_MUX_bit_math_h_l612_c3_b44b_cond,
layer0_node54_MUX_bit_math_h_l612_c3_b44b_iftrue,
layer0_node54_MUX_bit_math_h_l612_c3_b44b_iffalse,
layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output);

-- layer0_node55_MUX_bit_math_h_l623_c3_0aaf
layer0_node55_MUX_bit_math_h_l623_c3_0aaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node55_MUX_bit_math_h_l623_c3_0aaf_cond,
layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iftrue,
layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iffalse,
layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output);

-- layer0_node56_MUX_bit_math_h_l634_c3_6313
layer0_node56_MUX_bit_math_h_l634_c3_6313 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node56_MUX_bit_math_h_l634_c3_6313_cond,
layer0_node56_MUX_bit_math_h_l634_c3_6313_iftrue,
layer0_node56_MUX_bit_math_h_l634_c3_6313_iffalse,
layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output);

-- layer0_node57_MUX_bit_math_h_l645_c3_d8b1
layer0_node57_MUX_bit_math_h_l645_c3_d8b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node57_MUX_bit_math_h_l645_c3_d8b1_cond,
layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iftrue,
layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iffalse,
layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output);

-- layer0_node58_MUX_bit_math_h_l656_c3_485d
layer0_node58_MUX_bit_math_h_l656_c3_485d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node58_MUX_bit_math_h_l656_c3_485d_cond,
layer0_node58_MUX_bit_math_h_l656_c3_485d_iftrue,
layer0_node58_MUX_bit_math_h_l656_c3_485d_iffalse,
layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output);

-- layer0_node59_MUX_bit_math_h_l667_c3_6892
layer0_node59_MUX_bit_math_h_l667_c3_6892 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node59_MUX_bit_math_h_l667_c3_6892_cond,
layer0_node59_MUX_bit_math_h_l667_c3_6892_iftrue,
layer0_node59_MUX_bit_math_h_l667_c3_6892_iffalse,
layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output);

-- layer0_node60_MUX_bit_math_h_l678_c3_51ce
layer0_node60_MUX_bit_math_h_l678_c3_51ce : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node60_MUX_bit_math_h_l678_c3_51ce_cond,
layer0_node60_MUX_bit_math_h_l678_c3_51ce_iftrue,
layer0_node60_MUX_bit_math_h_l678_c3_51ce_iffalse,
layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output);

-- layer0_node61_MUX_bit_math_h_l689_c3_8d98
layer0_node61_MUX_bit_math_h_l689_c3_8d98 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node61_MUX_bit_math_h_l689_c3_8d98_cond,
layer0_node61_MUX_bit_math_h_l689_c3_8d98_iftrue,
layer0_node61_MUX_bit_math_h_l689_c3_8d98_iffalse,
layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output);

-- layer0_node62_MUX_bit_math_h_l700_c3_9327
layer0_node62_MUX_bit_math_h_l700_c3_9327 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node62_MUX_bit_math_h_l700_c3_9327_cond,
layer0_node62_MUX_bit_math_h_l700_c3_9327_iftrue,
layer0_node62_MUX_bit_math_h_l700_c3_9327_iffalse,
layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output);

-- layer0_node63_MUX_bit_math_h_l711_c3_c233
layer0_node63_MUX_bit_math_h_l711_c3_c233 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node63_MUX_bit_math_h_l711_c3_c233_cond,
layer0_node63_MUX_bit_math_h_l711_c3_c233_iftrue,
layer0_node63_MUX_bit_math_h_l711_c3_c233_iffalse,
layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output);

-- layer1_node0_MUX_bit_math_h_l728_c3_cd45
layer1_node0_MUX_bit_math_h_l728_c3_cd45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l728_c3_cd45_cond,
layer1_node0_MUX_bit_math_h_l728_c3_cd45_iftrue,
layer1_node0_MUX_bit_math_h_l728_c3_cd45_iffalse,
layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output);

-- layer1_node1_MUX_bit_math_h_l739_c3_e269
layer1_node1_MUX_bit_math_h_l739_c3_e269 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l739_c3_e269_cond,
layer1_node1_MUX_bit_math_h_l739_c3_e269_iftrue,
layer1_node1_MUX_bit_math_h_l739_c3_e269_iffalse,
layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output);

-- layer1_node2_MUX_bit_math_h_l750_c3_5aa6
layer1_node2_MUX_bit_math_h_l750_c3_5aa6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l750_c3_5aa6_cond,
layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iftrue,
layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iffalse,
layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output);

-- layer1_node3_MUX_bit_math_h_l761_c3_850a
layer1_node3_MUX_bit_math_h_l761_c3_850a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l761_c3_850a_cond,
layer1_node3_MUX_bit_math_h_l761_c3_850a_iftrue,
layer1_node3_MUX_bit_math_h_l761_c3_850a_iffalse,
layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output);

-- layer1_node4_MUX_bit_math_h_l772_c3_a071
layer1_node4_MUX_bit_math_h_l772_c3_a071 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node4_MUX_bit_math_h_l772_c3_a071_cond,
layer1_node4_MUX_bit_math_h_l772_c3_a071_iftrue,
layer1_node4_MUX_bit_math_h_l772_c3_a071_iffalse,
layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output);

-- layer1_node5_MUX_bit_math_h_l783_c3_9883
layer1_node5_MUX_bit_math_h_l783_c3_9883 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node5_MUX_bit_math_h_l783_c3_9883_cond,
layer1_node5_MUX_bit_math_h_l783_c3_9883_iftrue,
layer1_node5_MUX_bit_math_h_l783_c3_9883_iffalse,
layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output);

-- layer1_node6_MUX_bit_math_h_l794_c3_cf43
layer1_node6_MUX_bit_math_h_l794_c3_cf43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node6_MUX_bit_math_h_l794_c3_cf43_cond,
layer1_node6_MUX_bit_math_h_l794_c3_cf43_iftrue,
layer1_node6_MUX_bit_math_h_l794_c3_cf43_iffalse,
layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output);

-- layer1_node7_MUX_bit_math_h_l805_c3_c99c
layer1_node7_MUX_bit_math_h_l805_c3_c99c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node7_MUX_bit_math_h_l805_c3_c99c_cond,
layer1_node7_MUX_bit_math_h_l805_c3_c99c_iftrue,
layer1_node7_MUX_bit_math_h_l805_c3_c99c_iffalse,
layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output);

-- layer1_node8_MUX_bit_math_h_l816_c3_fa37
layer1_node8_MUX_bit_math_h_l816_c3_fa37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node8_MUX_bit_math_h_l816_c3_fa37_cond,
layer1_node8_MUX_bit_math_h_l816_c3_fa37_iftrue,
layer1_node8_MUX_bit_math_h_l816_c3_fa37_iffalse,
layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output);

-- layer1_node9_MUX_bit_math_h_l827_c3_d6c2
layer1_node9_MUX_bit_math_h_l827_c3_d6c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node9_MUX_bit_math_h_l827_c3_d6c2_cond,
layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iftrue,
layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iffalse,
layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output);

-- layer1_node10_MUX_bit_math_h_l838_c3_7eb8
layer1_node10_MUX_bit_math_h_l838_c3_7eb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node10_MUX_bit_math_h_l838_c3_7eb8_cond,
layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iftrue,
layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iffalse,
layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output);

-- layer1_node11_MUX_bit_math_h_l849_c3_2cb0
layer1_node11_MUX_bit_math_h_l849_c3_2cb0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node11_MUX_bit_math_h_l849_c3_2cb0_cond,
layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iftrue,
layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iffalse,
layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output);

-- layer1_node12_MUX_bit_math_h_l860_c3_32ef
layer1_node12_MUX_bit_math_h_l860_c3_32ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node12_MUX_bit_math_h_l860_c3_32ef_cond,
layer1_node12_MUX_bit_math_h_l860_c3_32ef_iftrue,
layer1_node12_MUX_bit_math_h_l860_c3_32ef_iffalse,
layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output);

-- layer1_node13_MUX_bit_math_h_l871_c3_c37d
layer1_node13_MUX_bit_math_h_l871_c3_c37d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node13_MUX_bit_math_h_l871_c3_c37d_cond,
layer1_node13_MUX_bit_math_h_l871_c3_c37d_iftrue,
layer1_node13_MUX_bit_math_h_l871_c3_c37d_iffalse,
layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output);

-- layer1_node14_MUX_bit_math_h_l882_c3_3e12
layer1_node14_MUX_bit_math_h_l882_c3_3e12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node14_MUX_bit_math_h_l882_c3_3e12_cond,
layer1_node14_MUX_bit_math_h_l882_c3_3e12_iftrue,
layer1_node14_MUX_bit_math_h_l882_c3_3e12_iffalse,
layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output);

-- layer1_node15_MUX_bit_math_h_l893_c3_5e2b
layer1_node15_MUX_bit_math_h_l893_c3_5e2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node15_MUX_bit_math_h_l893_c3_5e2b_cond,
layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iftrue,
layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iffalse,
layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output);

-- layer1_node16_MUX_bit_math_h_l904_c3_234e
layer1_node16_MUX_bit_math_h_l904_c3_234e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node16_MUX_bit_math_h_l904_c3_234e_cond,
layer1_node16_MUX_bit_math_h_l904_c3_234e_iftrue,
layer1_node16_MUX_bit_math_h_l904_c3_234e_iffalse,
layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output);

-- layer1_node17_MUX_bit_math_h_l915_c3_90a2
layer1_node17_MUX_bit_math_h_l915_c3_90a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node17_MUX_bit_math_h_l915_c3_90a2_cond,
layer1_node17_MUX_bit_math_h_l915_c3_90a2_iftrue,
layer1_node17_MUX_bit_math_h_l915_c3_90a2_iffalse,
layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output);

-- layer1_node18_MUX_bit_math_h_l926_c3_ecc8
layer1_node18_MUX_bit_math_h_l926_c3_ecc8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node18_MUX_bit_math_h_l926_c3_ecc8_cond,
layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iftrue,
layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iffalse,
layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output);

-- layer1_node19_MUX_bit_math_h_l937_c3_7211
layer1_node19_MUX_bit_math_h_l937_c3_7211 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node19_MUX_bit_math_h_l937_c3_7211_cond,
layer1_node19_MUX_bit_math_h_l937_c3_7211_iftrue,
layer1_node19_MUX_bit_math_h_l937_c3_7211_iffalse,
layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output);

-- layer1_node20_MUX_bit_math_h_l948_c3_2d00
layer1_node20_MUX_bit_math_h_l948_c3_2d00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node20_MUX_bit_math_h_l948_c3_2d00_cond,
layer1_node20_MUX_bit_math_h_l948_c3_2d00_iftrue,
layer1_node20_MUX_bit_math_h_l948_c3_2d00_iffalse,
layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output);

-- layer1_node21_MUX_bit_math_h_l959_c3_f682
layer1_node21_MUX_bit_math_h_l959_c3_f682 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node21_MUX_bit_math_h_l959_c3_f682_cond,
layer1_node21_MUX_bit_math_h_l959_c3_f682_iftrue,
layer1_node21_MUX_bit_math_h_l959_c3_f682_iffalse,
layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output);

-- layer1_node22_MUX_bit_math_h_l970_c3_8998
layer1_node22_MUX_bit_math_h_l970_c3_8998 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node22_MUX_bit_math_h_l970_c3_8998_cond,
layer1_node22_MUX_bit_math_h_l970_c3_8998_iftrue,
layer1_node22_MUX_bit_math_h_l970_c3_8998_iffalse,
layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output);

-- layer1_node23_MUX_bit_math_h_l981_c3_102a
layer1_node23_MUX_bit_math_h_l981_c3_102a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node23_MUX_bit_math_h_l981_c3_102a_cond,
layer1_node23_MUX_bit_math_h_l981_c3_102a_iftrue,
layer1_node23_MUX_bit_math_h_l981_c3_102a_iffalse,
layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output);

-- layer1_node24_MUX_bit_math_h_l992_c3_9fd6
layer1_node24_MUX_bit_math_h_l992_c3_9fd6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node24_MUX_bit_math_h_l992_c3_9fd6_cond,
layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iftrue,
layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iffalse,
layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output);

-- layer1_node25_MUX_bit_math_h_l1003_c3_271e
layer1_node25_MUX_bit_math_h_l1003_c3_271e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node25_MUX_bit_math_h_l1003_c3_271e_cond,
layer1_node25_MUX_bit_math_h_l1003_c3_271e_iftrue,
layer1_node25_MUX_bit_math_h_l1003_c3_271e_iffalse,
layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output);

-- layer1_node26_MUX_bit_math_h_l1014_c3_1e7d
layer1_node26_MUX_bit_math_h_l1014_c3_1e7d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_cond,
layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iftrue,
layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iffalse,
layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output);

-- layer1_node27_MUX_bit_math_h_l1025_c3_46dd
layer1_node27_MUX_bit_math_h_l1025_c3_46dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node27_MUX_bit_math_h_l1025_c3_46dd_cond,
layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iftrue,
layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iffalse,
layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output);

-- layer1_node28_MUX_bit_math_h_l1036_c3_4035
layer1_node28_MUX_bit_math_h_l1036_c3_4035 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node28_MUX_bit_math_h_l1036_c3_4035_cond,
layer1_node28_MUX_bit_math_h_l1036_c3_4035_iftrue,
layer1_node28_MUX_bit_math_h_l1036_c3_4035_iffalse,
layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output);

-- layer1_node29_MUX_bit_math_h_l1047_c3_3314
layer1_node29_MUX_bit_math_h_l1047_c3_3314 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node29_MUX_bit_math_h_l1047_c3_3314_cond,
layer1_node29_MUX_bit_math_h_l1047_c3_3314_iftrue,
layer1_node29_MUX_bit_math_h_l1047_c3_3314_iffalse,
layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output);

-- layer1_node30_MUX_bit_math_h_l1058_c3_6a5f
layer1_node30_MUX_bit_math_h_l1058_c3_6a5f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_cond,
layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iftrue,
layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iffalse,
layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output);

-- layer1_node31_MUX_bit_math_h_l1069_c3_5488
layer1_node31_MUX_bit_math_h_l1069_c3_5488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node31_MUX_bit_math_h_l1069_c3_5488_cond,
layer1_node31_MUX_bit_math_h_l1069_c3_5488_iftrue,
layer1_node31_MUX_bit_math_h_l1069_c3_5488_iffalse,
layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output);

-- layer2_node0_MUX_bit_math_h_l1086_c3_74df
layer2_node0_MUX_bit_math_h_l1086_c3_74df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l1086_c3_74df_cond,
layer2_node0_MUX_bit_math_h_l1086_c3_74df_iftrue,
layer2_node0_MUX_bit_math_h_l1086_c3_74df_iffalse,
layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output);

-- layer2_node1_MUX_bit_math_h_l1097_c3_4739
layer2_node1_MUX_bit_math_h_l1097_c3_4739 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l1097_c3_4739_cond,
layer2_node1_MUX_bit_math_h_l1097_c3_4739_iftrue,
layer2_node1_MUX_bit_math_h_l1097_c3_4739_iffalse,
layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output);

-- layer2_node2_MUX_bit_math_h_l1108_c3_c83e
layer2_node2_MUX_bit_math_h_l1108_c3_c83e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node2_MUX_bit_math_h_l1108_c3_c83e_cond,
layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iftrue,
layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iffalse,
layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output);

-- layer2_node3_MUX_bit_math_h_l1119_c3_1d4a
layer2_node3_MUX_bit_math_h_l1119_c3_1d4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_cond,
layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iftrue,
layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iffalse,
layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output);

-- layer2_node4_MUX_bit_math_h_l1130_c3_d0b7
layer2_node4_MUX_bit_math_h_l1130_c3_d0b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_cond,
layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iftrue,
layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iffalse,
layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output);

-- layer2_node5_MUX_bit_math_h_l1141_c3_a33d
layer2_node5_MUX_bit_math_h_l1141_c3_a33d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node5_MUX_bit_math_h_l1141_c3_a33d_cond,
layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iftrue,
layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iffalse,
layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output);

-- layer2_node6_MUX_bit_math_h_l1152_c3_403d
layer2_node6_MUX_bit_math_h_l1152_c3_403d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node6_MUX_bit_math_h_l1152_c3_403d_cond,
layer2_node6_MUX_bit_math_h_l1152_c3_403d_iftrue,
layer2_node6_MUX_bit_math_h_l1152_c3_403d_iffalse,
layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output);

-- layer2_node7_MUX_bit_math_h_l1163_c3_f8a3
layer2_node7_MUX_bit_math_h_l1163_c3_f8a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_cond,
layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iftrue,
layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iffalse,
layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output);

-- layer2_node8_MUX_bit_math_h_l1174_c3_51d4
layer2_node8_MUX_bit_math_h_l1174_c3_51d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node8_MUX_bit_math_h_l1174_c3_51d4_cond,
layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iftrue,
layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iffalse,
layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output);

-- layer2_node9_MUX_bit_math_h_l1185_c3_30b5
layer2_node9_MUX_bit_math_h_l1185_c3_30b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node9_MUX_bit_math_h_l1185_c3_30b5_cond,
layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iftrue,
layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iffalse,
layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output);

-- layer2_node10_MUX_bit_math_h_l1196_c3_6142
layer2_node10_MUX_bit_math_h_l1196_c3_6142 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node10_MUX_bit_math_h_l1196_c3_6142_cond,
layer2_node10_MUX_bit_math_h_l1196_c3_6142_iftrue,
layer2_node10_MUX_bit_math_h_l1196_c3_6142_iffalse,
layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output);

-- layer2_node11_MUX_bit_math_h_l1207_c3_17d4
layer2_node11_MUX_bit_math_h_l1207_c3_17d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node11_MUX_bit_math_h_l1207_c3_17d4_cond,
layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iftrue,
layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iffalse,
layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output);

-- layer2_node12_MUX_bit_math_h_l1218_c3_74f5
layer2_node12_MUX_bit_math_h_l1218_c3_74f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node12_MUX_bit_math_h_l1218_c3_74f5_cond,
layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iftrue,
layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iffalse,
layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output);

-- layer2_node13_MUX_bit_math_h_l1229_c3_af85
layer2_node13_MUX_bit_math_h_l1229_c3_af85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node13_MUX_bit_math_h_l1229_c3_af85_cond,
layer2_node13_MUX_bit_math_h_l1229_c3_af85_iftrue,
layer2_node13_MUX_bit_math_h_l1229_c3_af85_iffalse,
layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output);

-- layer2_node14_MUX_bit_math_h_l1240_c3_0287
layer2_node14_MUX_bit_math_h_l1240_c3_0287 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node14_MUX_bit_math_h_l1240_c3_0287_cond,
layer2_node14_MUX_bit_math_h_l1240_c3_0287_iftrue,
layer2_node14_MUX_bit_math_h_l1240_c3_0287_iffalse,
layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output);

-- layer2_node15_MUX_bit_math_h_l1251_c3_a113
layer2_node15_MUX_bit_math_h_l1251_c3_a113 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node15_MUX_bit_math_h_l1251_c3_a113_cond,
layer2_node15_MUX_bit_math_h_l1251_c3_a113_iftrue,
layer2_node15_MUX_bit_math_h_l1251_c3_a113_iffalse,
layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output);

-- layer3_node0_MUX_bit_math_h_l1268_c3_1d33
layer3_node0_MUX_bit_math_h_l1268_c3_1d33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l1268_c3_1d33_cond,
layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iftrue,
layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iffalse,
layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output);

-- layer3_node1_MUX_bit_math_h_l1279_c3_ca08
layer3_node1_MUX_bit_math_h_l1279_c3_ca08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node1_MUX_bit_math_h_l1279_c3_ca08_cond,
layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iftrue,
layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iffalse,
layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output);

-- layer3_node2_MUX_bit_math_h_l1290_c3_581b
layer3_node2_MUX_bit_math_h_l1290_c3_581b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node2_MUX_bit_math_h_l1290_c3_581b_cond,
layer3_node2_MUX_bit_math_h_l1290_c3_581b_iftrue,
layer3_node2_MUX_bit_math_h_l1290_c3_581b_iffalse,
layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output);

-- layer3_node3_MUX_bit_math_h_l1301_c3_778a
layer3_node3_MUX_bit_math_h_l1301_c3_778a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node3_MUX_bit_math_h_l1301_c3_778a_cond,
layer3_node3_MUX_bit_math_h_l1301_c3_778a_iftrue,
layer3_node3_MUX_bit_math_h_l1301_c3_778a_iffalse,
layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output);

-- layer3_node4_MUX_bit_math_h_l1312_c3_9af8
layer3_node4_MUX_bit_math_h_l1312_c3_9af8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node4_MUX_bit_math_h_l1312_c3_9af8_cond,
layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iftrue,
layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iffalse,
layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output);

-- layer3_node5_MUX_bit_math_h_l1323_c3_8487
layer3_node5_MUX_bit_math_h_l1323_c3_8487 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node5_MUX_bit_math_h_l1323_c3_8487_cond,
layer3_node5_MUX_bit_math_h_l1323_c3_8487_iftrue,
layer3_node5_MUX_bit_math_h_l1323_c3_8487_iffalse,
layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output);

-- layer3_node6_MUX_bit_math_h_l1334_c3_d703
layer3_node6_MUX_bit_math_h_l1334_c3_d703 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node6_MUX_bit_math_h_l1334_c3_d703_cond,
layer3_node6_MUX_bit_math_h_l1334_c3_d703_iftrue,
layer3_node6_MUX_bit_math_h_l1334_c3_d703_iffalse,
layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output);

-- layer3_node7_MUX_bit_math_h_l1345_c3_ae83
layer3_node7_MUX_bit_math_h_l1345_c3_ae83 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node7_MUX_bit_math_h_l1345_c3_ae83_cond,
layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iftrue,
layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iffalse,
layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output);

-- layer4_node0_MUX_bit_math_h_l1362_c3_0390
layer4_node0_MUX_bit_math_h_l1362_c3_0390 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node0_MUX_bit_math_h_l1362_c3_0390_cond,
layer4_node0_MUX_bit_math_h_l1362_c3_0390_iftrue,
layer4_node0_MUX_bit_math_h_l1362_c3_0390_iffalse,
layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output);

-- layer4_node1_MUX_bit_math_h_l1373_c3_27d5
layer4_node1_MUX_bit_math_h_l1373_c3_27d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node1_MUX_bit_math_h_l1373_c3_27d5_cond,
layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iftrue,
layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iffalse,
layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output);

-- layer4_node2_MUX_bit_math_h_l1384_c3_2032
layer4_node2_MUX_bit_math_h_l1384_c3_2032 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node2_MUX_bit_math_h_l1384_c3_2032_cond,
layer4_node2_MUX_bit_math_h_l1384_c3_2032_iftrue,
layer4_node2_MUX_bit_math_h_l1384_c3_2032_iffalse,
layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output);

-- layer4_node3_MUX_bit_math_h_l1395_c3_ef44
layer4_node3_MUX_bit_math_h_l1395_c3_ef44 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node3_MUX_bit_math_h_l1395_c3_ef44_cond,
layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iftrue,
layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iffalse,
layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output);

-- layer5_node0_MUX_bit_math_h_l1412_c3_1733
layer5_node0_MUX_bit_math_h_l1412_c3_1733 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node0_MUX_bit_math_h_l1412_c3_1733_cond,
layer5_node0_MUX_bit_math_h_l1412_c3_1733_iftrue,
layer5_node0_MUX_bit_math_h_l1412_c3_1733_iffalse,
layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output);

-- layer5_node1_MUX_bit_math_h_l1423_c3_54e8
layer5_node1_MUX_bit_math_h_l1423_c3_54e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node1_MUX_bit_math_h_l1423_c3_54e8_cond,
layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iftrue,
layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iffalse,
layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output);

-- layer6_node0_MUX_bit_math_h_l1440_c3_c11f
layer6_node0_MUX_bit_math_h_l1440_c3_c11f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer6_node0_MUX_bit_math_h_l1440_c3_c11f_cond,
layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iftrue,
layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iffalse,
layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 in16,
 in17,
 in18,
 in19,
 in20,
 in21,
 in22,
 in23,
 in24,
 in25,
 in26,
 in27,
 in28,
 in29,
 in30,
 in31,
 in32,
 in33,
 in34,
 in35,
 in36,
 in37,
 in38,
 in39,
 in40,
 in41,
 in42,
 in43,
 in44,
 in45,
 in46,
 in47,
 in48,
 in49,
 in50,
 in51,
 in52,
 in53,
 in54,
 in55,
 in56,
 in57,
 in58,
 in59,
 in60,
 in61,
 in62,
 in63,
 in64,
 in65,
 in66,
 in67,
 in68,
 in69,
 in70,
 in71,
 in72,
 in73,
 in74,
 in75,
 in76,
 in77,
 in78,
 in79,
 in80,
 in81,
 in82,
 in83,
 in84,
 in85,
 in86,
 in87,
 in88,
 in89,
 in90,
 in91,
 in92,
 in93,
 in94,
 in95,
 in96,
 in97,
 in98,
 in99,
 in100,
 in101,
 in102,
 in103,
 in104,
 in105,
 in106,
 in107,
 in108,
 in109,
 in110,
 in111,
 in112,
 in113,
 in114,
 in115,
 in116,
 in117,
 in118,
 in119,
 in120,
 in121,
 in122,
 in123,
 in124,
 in125,
 in126,
 in127,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output,
 layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output,
 layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output,
 layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output,
 layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output,
 layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output,
 layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output,
 layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output,
 layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output,
 layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output,
 layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output,
 layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output,
 layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output,
 layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output,
 layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output,
 layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output,
 layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output,
 layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output,
 layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output,
 layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output,
 layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output,
 layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output,
 layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output,
 layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output,
 layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output,
 layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output,
 layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output,
 layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output,
 layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output,
 layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output,
 layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output,
 layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output,
 layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output,
 layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output,
 layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output,
 layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output,
 layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output,
 layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output,
 layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output,
 layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output,
 layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output,
 layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output,
 layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output,
 layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output,
 layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output,
 layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output,
 layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output,
 layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output,
 layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output,
 layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output,
 layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output,
 layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output,
 layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output,
 layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output,
 layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output,
 layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output,
 layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output,
 layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output,
 layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output,
 layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output,
 layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output,
 layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output,
 layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output,
 layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output,
 layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output,
 layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output,
 layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output,
 layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output,
 layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output,
 layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output,
 layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output,
 layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output,
 layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output,
 layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output,
 layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output,
 layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output,
 layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output,
 layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output,
 layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output,
 layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output,
 layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output,
 layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output,
 layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output,
 layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output,
 layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output,
 layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output,
 layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output,
 layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output,
 layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output,
 layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output,
 layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output,
 layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output,
 layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output,
 layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output,
 layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output,
 layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output,
 layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output,
 layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output,
 layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output,
 layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output,
 layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output,
 layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output,
 layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output,
 layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output,
 layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output,
 layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output,
 layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output,
 layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output,
 layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output,
 layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output,
 layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output,
 layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output,
 layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output,
 layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output,
 layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output,
 layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output,
 layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output,
 layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output,
 layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output,
 layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_in0 : unsigned(7 downto 0);
 variable VAR_in1 : unsigned(7 downto 0);
 variable VAR_in2 : unsigned(7 downto 0);
 variable VAR_in3 : unsigned(7 downto 0);
 variable VAR_in4 : unsigned(7 downto 0);
 variable VAR_in5 : unsigned(7 downto 0);
 variable VAR_in6 : unsigned(7 downto 0);
 variable VAR_in7 : unsigned(7 downto 0);
 variable VAR_in8 : unsigned(7 downto 0);
 variable VAR_in9 : unsigned(7 downto 0);
 variable VAR_in10 : unsigned(7 downto 0);
 variable VAR_in11 : unsigned(7 downto 0);
 variable VAR_in12 : unsigned(7 downto 0);
 variable VAR_in13 : unsigned(7 downto 0);
 variable VAR_in14 : unsigned(7 downto 0);
 variable VAR_in15 : unsigned(7 downto 0);
 variable VAR_in16 : unsigned(7 downto 0);
 variable VAR_in17 : unsigned(7 downto 0);
 variable VAR_in18 : unsigned(7 downto 0);
 variable VAR_in19 : unsigned(7 downto 0);
 variable VAR_in20 : unsigned(7 downto 0);
 variable VAR_in21 : unsigned(7 downto 0);
 variable VAR_in22 : unsigned(7 downto 0);
 variable VAR_in23 : unsigned(7 downto 0);
 variable VAR_in24 : unsigned(7 downto 0);
 variable VAR_in25 : unsigned(7 downto 0);
 variable VAR_in26 : unsigned(7 downto 0);
 variable VAR_in27 : unsigned(7 downto 0);
 variable VAR_in28 : unsigned(7 downto 0);
 variable VAR_in29 : unsigned(7 downto 0);
 variable VAR_in30 : unsigned(7 downto 0);
 variable VAR_in31 : unsigned(7 downto 0);
 variable VAR_in32 : unsigned(7 downto 0);
 variable VAR_in33 : unsigned(7 downto 0);
 variable VAR_in34 : unsigned(7 downto 0);
 variable VAR_in35 : unsigned(7 downto 0);
 variable VAR_in36 : unsigned(7 downto 0);
 variable VAR_in37 : unsigned(7 downto 0);
 variable VAR_in38 : unsigned(7 downto 0);
 variable VAR_in39 : unsigned(7 downto 0);
 variable VAR_in40 : unsigned(7 downto 0);
 variable VAR_in41 : unsigned(7 downto 0);
 variable VAR_in42 : unsigned(7 downto 0);
 variable VAR_in43 : unsigned(7 downto 0);
 variable VAR_in44 : unsigned(7 downto 0);
 variable VAR_in45 : unsigned(7 downto 0);
 variable VAR_in46 : unsigned(7 downto 0);
 variable VAR_in47 : unsigned(7 downto 0);
 variable VAR_in48 : unsigned(7 downto 0);
 variable VAR_in49 : unsigned(7 downto 0);
 variable VAR_in50 : unsigned(7 downto 0);
 variable VAR_in51 : unsigned(7 downto 0);
 variable VAR_in52 : unsigned(7 downto 0);
 variable VAR_in53 : unsigned(7 downto 0);
 variable VAR_in54 : unsigned(7 downto 0);
 variable VAR_in55 : unsigned(7 downto 0);
 variable VAR_in56 : unsigned(7 downto 0);
 variable VAR_in57 : unsigned(7 downto 0);
 variable VAR_in58 : unsigned(7 downto 0);
 variable VAR_in59 : unsigned(7 downto 0);
 variable VAR_in60 : unsigned(7 downto 0);
 variable VAR_in61 : unsigned(7 downto 0);
 variable VAR_in62 : unsigned(7 downto 0);
 variable VAR_in63 : unsigned(7 downto 0);
 variable VAR_in64 : unsigned(7 downto 0);
 variable VAR_in65 : unsigned(7 downto 0);
 variable VAR_in66 : unsigned(7 downto 0);
 variable VAR_in67 : unsigned(7 downto 0);
 variable VAR_in68 : unsigned(7 downto 0);
 variable VAR_in69 : unsigned(7 downto 0);
 variable VAR_in70 : unsigned(7 downto 0);
 variable VAR_in71 : unsigned(7 downto 0);
 variable VAR_in72 : unsigned(7 downto 0);
 variable VAR_in73 : unsigned(7 downto 0);
 variable VAR_in74 : unsigned(7 downto 0);
 variable VAR_in75 : unsigned(7 downto 0);
 variable VAR_in76 : unsigned(7 downto 0);
 variable VAR_in77 : unsigned(7 downto 0);
 variable VAR_in78 : unsigned(7 downto 0);
 variable VAR_in79 : unsigned(7 downto 0);
 variable VAR_in80 : unsigned(7 downto 0);
 variable VAR_in81 : unsigned(7 downto 0);
 variable VAR_in82 : unsigned(7 downto 0);
 variable VAR_in83 : unsigned(7 downto 0);
 variable VAR_in84 : unsigned(7 downto 0);
 variable VAR_in85 : unsigned(7 downto 0);
 variable VAR_in86 : unsigned(7 downto 0);
 variable VAR_in87 : unsigned(7 downto 0);
 variable VAR_in88 : unsigned(7 downto 0);
 variable VAR_in89 : unsigned(7 downto 0);
 variable VAR_in90 : unsigned(7 downto 0);
 variable VAR_in91 : unsigned(7 downto 0);
 variable VAR_in92 : unsigned(7 downto 0);
 variable VAR_in93 : unsigned(7 downto 0);
 variable VAR_in94 : unsigned(7 downto 0);
 variable VAR_in95 : unsigned(7 downto 0);
 variable VAR_in96 : unsigned(7 downto 0);
 variable VAR_in97 : unsigned(7 downto 0);
 variable VAR_in98 : unsigned(7 downto 0);
 variable VAR_in99 : unsigned(7 downto 0);
 variable VAR_in100 : unsigned(7 downto 0);
 variable VAR_in101 : unsigned(7 downto 0);
 variable VAR_in102 : unsigned(7 downto 0);
 variable VAR_in103 : unsigned(7 downto 0);
 variable VAR_in104 : unsigned(7 downto 0);
 variable VAR_in105 : unsigned(7 downto 0);
 variable VAR_in106 : unsigned(7 downto 0);
 variable VAR_in107 : unsigned(7 downto 0);
 variable VAR_in108 : unsigned(7 downto 0);
 variable VAR_in109 : unsigned(7 downto 0);
 variable VAR_in110 : unsigned(7 downto 0);
 variable VAR_in111 : unsigned(7 downto 0);
 variable VAR_in112 : unsigned(7 downto 0);
 variable VAR_in113 : unsigned(7 downto 0);
 variable VAR_in114 : unsigned(7 downto 0);
 variable VAR_in115 : unsigned(7 downto 0);
 variable VAR_in116 : unsigned(7 downto 0);
 variable VAR_in117 : unsigned(7 downto 0);
 variable VAR_in118 : unsigned(7 downto 0);
 variable VAR_in119 : unsigned(7 downto 0);
 variable VAR_in120 : unsigned(7 downto 0);
 variable VAR_in121 : unsigned(7 downto 0);
 variable VAR_in122 : unsigned(7 downto 0);
 variable VAR_in123 : unsigned(7 downto 0);
 variable VAR_in124 : unsigned(7 downto 0);
 variable VAR_in125 : unsigned(7 downto 0);
 variable VAR_in126 : unsigned(7 downto 0);
 variable VAR_in127 : unsigned(7 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_cond : unsigned(0 downto 0);
 variable VAR_layer0_node8 : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_cond : unsigned(0 downto 0);
 variable VAR_layer0_node9 : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node10 : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_cond : unsigned(0 downto 0);
 variable VAR_layer0_node11 : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node12 : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_cond : unsigned(0 downto 0);
 variable VAR_layer0_node13 : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node14 : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_cond : unsigned(0 downto 0);
 variable VAR_layer0_node15 : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_cond : unsigned(0 downto 0);
 variable VAR_layer0_node16 : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_cond : unsigned(0 downto 0);
 variable VAR_layer0_node17 : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node18 : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_cond : unsigned(0 downto 0);
 variable VAR_layer0_node19 : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_cond : unsigned(0 downto 0);
 variable VAR_layer0_node20 : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node21 : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_cond : unsigned(0 downto 0);
 variable VAR_layer0_node22 : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_cond : unsigned(0 downto 0);
 variable VAR_layer0_node23 : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node24 : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_cond : unsigned(0 downto 0);
 variable VAR_layer0_node25 : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node26 : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node27 : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node28 : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_cond : unsigned(0 downto 0);
 variable VAR_layer0_node29 : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_cond : unsigned(0 downto 0);
 variable VAR_layer0_node30 : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_cond : unsigned(0 downto 0);
 variable VAR_layer0_node31 : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_cond : unsigned(0 downto 0);
 variable VAR_layer0_node32 : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_cond : unsigned(0 downto 0);
 variable VAR_layer0_node33 : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_cond : unsigned(0 downto 0);
 variable VAR_layer0_node34 : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_cond : unsigned(0 downto 0);
 variable VAR_layer0_node35 : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node36 : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_cond : unsigned(0 downto 0);
 variable VAR_layer0_node37 : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_cond : unsigned(0 downto 0);
 variable VAR_layer0_node38 : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_cond : unsigned(0 downto 0);
 variable VAR_layer0_node39 : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node40 : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_cond : unsigned(0 downto 0);
 variable VAR_layer0_node41 : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_cond : unsigned(0 downto 0);
 variable VAR_layer0_node42 : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node43 : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_cond : unsigned(0 downto 0);
 variable VAR_layer0_node44 : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node45 : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node46 : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_cond : unsigned(0 downto 0);
 variable VAR_layer0_node47 : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_cond : unsigned(0 downto 0);
 variable VAR_layer0_node48 : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_cond : unsigned(0 downto 0);
 variable VAR_layer0_node49 : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node50 : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_cond : unsigned(0 downto 0);
 variable VAR_layer0_node51 : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node52 : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node53 : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node54 : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node55 : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_cond : unsigned(0 downto 0);
 variable VAR_layer0_node56 : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_cond : unsigned(0 downto 0);
 variable VAR_layer0_node57 : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node58 : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node59 : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_cond : unsigned(0 downto 0);
 variable VAR_layer0_node60 : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_cond : unsigned(0 downto 0);
 variable VAR_layer0_node61 : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_cond : unsigned(0 downto 0);
 variable VAR_layer0_node62 : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_cond : unsigned(0 downto 0);
 variable VAR_layer0_node63 : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node4 : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_cond : unsigned(0 downto 0);
 variable VAR_layer1_node5 : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_cond : unsigned(0 downto 0);
 variable VAR_layer1_node6 : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_cond : unsigned(0 downto 0);
 variable VAR_layer1_node7 : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_cond : unsigned(0 downto 0);
 variable VAR_layer1_node8 : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_cond : unsigned(0 downto 0);
 variable VAR_layer1_node9 : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_cond : unsigned(0 downto 0);
 variable VAR_layer1_node10 : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_cond : unsigned(0 downto 0);
 variable VAR_layer1_node11 : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_cond : unsigned(0 downto 0);
 variable VAR_layer1_node12 : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_cond : unsigned(0 downto 0);
 variable VAR_layer1_node13 : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node14 : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_cond : unsigned(0 downto 0);
 variable VAR_layer1_node15 : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_cond : unsigned(0 downto 0);
 variable VAR_layer1_node16 : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_cond : unsigned(0 downto 0);
 variable VAR_layer1_node17 : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_cond : unsigned(0 downto 0);
 variable VAR_layer1_node18 : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_cond : unsigned(0 downto 0);
 variable VAR_layer1_node19 : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_cond : unsigned(0 downto 0);
 variable VAR_layer1_node20 : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_cond : unsigned(0 downto 0);
 variable VAR_layer1_node21 : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_cond : unsigned(0 downto 0);
 variable VAR_layer1_node22 : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_cond : unsigned(0 downto 0);
 variable VAR_layer1_node23 : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node24 : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_cond : unsigned(0 downto 0);
 variable VAR_layer1_node25 : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_cond : unsigned(0 downto 0);
 variable VAR_layer1_node26 : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node27 : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_cond : unsigned(0 downto 0);
 variable VAR_layer1_node28 : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_cond : unsigned(0 downto 0);
 variable VAR_layer1_node29 : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_cond : unsigned(0 downto 0);
 variable VAR_layer1_node30 : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node31 : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_cond : unsigned(0 downto 0);
 variable VAR_layer2_node2 : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_cond : unsigned(0 downto 0);
 variable VAR_layer2_node3 : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_cond : unsigned(0 downto 0);
 variable VAR_layer2_node4 : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_cond : unsigned(0 downto 0);
 variable VAR_layer2_node5 : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node6 : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node7 : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_cond : unsigned(0 downto 0);
 variable VAR_layer2_node8 : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_cond : unsigned(0 downto 0);
 variable VAR_layer2_node9 : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_cond : unsigned(0 downto 0);
 variable VAR_layer2_node10 : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_cond : unsigned(0 downto 0);
 variable VAR_layer2_node11 : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_cond : unsigned(0 downto 0);
 variable VAR_layer2_node12 : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_cond : unsigned(0 downto 0);
 variable VAR_layer2_node13 : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_cond : unsigned(0 downto 0);
 variable VAR_layer2_node14 : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_cond : unsigned(0 downto 0);
 variable VAR_layer2_node15 : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_cond : unsigned(0 downto 0);
 variable VAR_layer3_node1 : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_cond : unsigned(0 downto 0);
 variable VAR_layer3_node2 : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_cond : unsigned(0 downto 0);
 variable VAR_layer3_node3 : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_cond : unsigned(0 downto 0);
 variable VAR_layer3_node4 : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_cond : unsigned(0 downto 0);
 variable VAR_layer3_node5 : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_cond : unsigned(0 downto 0);
 variable VAR_layer3_node6 : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_cond : unsigned(0 downto 0);
 variable VAR_layer3_node7 : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_cond : unsigned(0 downto 0);
 variable VAR_sel4 : unsigned(0 downto 0);
 variable VAR_uint7_4_4_bit_math_h_l1358_c10_39f5_return_output : unsigned(0 downto 0);
 variable VAR_layer4_node0 : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_cond : unsigned(0 downto 0);
 variable VAR_layer4_node1 : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_cond : unsigned(0 downto 0);
 variable VAR_layer4_node2 : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_cond : unsigned(0 downto 0);
 variable VAR_layer4_node3 : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_cond : unsigned(0 downto 0);
 variable VAR_sel5 : unsigned(0 downto 0);
 variable VAR_uint7_5_5_bit_math_h_l1408_c10_5487_return_output : unsigned(0 downto 0);
 variable VAR_layer5_node0 : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_cond : unsigned(0 downto 0);
 variable VAR_layer5_node1 : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_cond : unsigned(0 downto 0);
 variable VAR_sel6 : unsigned(0 downto 0);
 variable VAR_uint7_6_6_bit_math_h_l1436_c10_41fb_return_output : unsigned(0 downto 0);
 variable VAR_layer6_node0 : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iftrue : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iffalse : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;
     VAR_in16 := in16;
     VAR_in17 := in17;
     VAR_in18 := in18;
     VAR_in19 := in19;
     VAR_in20 := in20;
     VAR_in21 := in21;
     VAR_in22 := in22;
     VAR_in23 := in23;
     VAR_in24 := in24;
     VAR_in25 := in25;
     VAR_in26 := in26;
     VAR_in27 := in27;
     VAR_in28 := in28;
     VAR_in29 := in29;
     VAR_in30 := in30;
     VAR_in31 := in31;
     VAR_in32 := in32;
     VAR_in33 := in33;
     VAR_in34 := in34;
     VAR_in35 := in35;
     VAR_in36 := in36;
     VAR_in37 := in37;
     VAR_in38 := in38;
     VAR_in39 := in39;
     VAR_in40 := in40;
     VAR_in41 := in41;
     VAR_in42 := in42;
     VAR_in43 := in43;
     VAR_in44 := in44;
     VAR_in45 := in45;
     VAR_in46 := in46;
     VAR_in47 := in47;
     VAR_in48 := in48;
     VAR_in49 := in49;
     VAR_in50 := in50;
     VAR_in51 := in51;
     VAR_in52 := in52;
     VAR_in53 := in53;
     VAR_in54 := in54;
     VAR_in55 := in55;
     VAR_in56 := in56;
     VAR_in57 := in57;
     VAR_in58 := in58;
     VAR_in59 := in59;
     VAR_in60 := in60;
     VAR_in61 := in61;
     VAR_in62 := in62;
     VAR_in63 := in63;
     VAR_in64 := in64;
     VAR_in65 := in65;
     VAR_in66 := in66;
     VAR_in67 := in67;
     VAR_in68 := in68;
     VAR_in69 := in69;
     VAR_in70 := in70;
     VAR_in71 := in71;
     VAR_in72 := in72;
     VAR_in73 := in73;
     VAR_in74 := in74;
     VAR_in75 := in75;
     VAR_in76 := in76;
     VAR_in77 := in77;
     VAR_in78 := in78;
     VAR_in79 := in79;
     VAR_in80 := in80;
     VAR_in81 := in81;
     VAR_in82 := in82;
     VAR_in83 := in83;
     VAR_in84 := in84;
     VAR_in85 := in85;
     VAR_in86 := in86;
     VAR_in87 := in87;
     VAR_in88 := in88;
     VAR_in89 := in89;
     VAR_in90 := in90;
     VAR_in91 := in91;
     VAR_in92 := in92;
     VAR_in93 := in93;
     VAR_in94 := in94;
     VAR_in95 := in95;
     VAR_in96 := in96;
     VAR_in97 := in97;
     VAR_in98 := in98;
     VAR_in99 := in99;
     VAR_in100 := in100;
     VAR_in101 := in101;
     VAR_in102 := in102;
     VAR_in103 := in103;
     VAR_in104 := in104;
     VAR_in105 := in105;
     VAR_in106 := in106;
     VAR_in107 := in107;
     VAR_in108 := in108;
     VAR_in109 := in109;
     VAR_in110 := in110;
     VAR_in111 := in111;
     VAR_in112 := in112;
     VAR_in113 := in113;
     VAR_in114 := in114;
     VAR_in115 := in115;
     VAR_in116 := in116;
     VAR_in117 := in117;
     VAR_in118 := in118;
     VAR_in119 := in119;
     VAR_in120 := in120;
     VAR_in121 := in121;
     VAR_in122 := in122;
     VAR_in123 := in123;
     VAR_in124 := in124;
     VAR_in125 := in125;
     VAR_in126 := in126;
     VAR_in127 := in127;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iffalse := VAR_in10;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_iffalse := VAR_in100;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_iftrue := VAR_in101;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_iffalse := VAR_in102;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_iftrue := VAR_in103;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iffalse := VAR_in104;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iftrue := VAR_in105;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_iffalse := VAR_in106;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_iftrue := VAR_in107;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_iffalse := VAR_in108;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_iftrue := VAR_in109;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iftrue := VAR_in11;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iffalse := VAR_in110;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iftrue := VAR_in111;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_iffalse := VAR_in112;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_iftrue := VAR_in113;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iffalse := VAR_in114;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iftrue := VAR_in115;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_iffalse := VAR_in116;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_iftrue := VAR_in117;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_iffalse := VAR_in118;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_iftrue := VAR_in119;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_iffalse := VAR_in12;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_iffalse := VAR_in120;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_iftrue := VAR_in121;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_iffalse := VAR_in122;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_iftrue := VAR_in123;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_iffalse := VAR_in124;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_iftrue := VAR_in125;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_iffalse := VAR_in126;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_iftrue := VAR_in127;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_iftrue := VAR_in15;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_iffalse := VAR_in16;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_iftrue := VAR_in17;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_iffalse := VAR_in18;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_iftrue := VAR_in19;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_iffalse := VAR_in2;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_iffalse := VAR_in20;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_iftrue := VAR_in21;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_iffalse := VAR_in22;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_iftrue := VAR_in23;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_iffalse := VAR_in24;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_iftrue := VAR_in25;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_iffalse := VAR_in26;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_iftrue := VAR_in27;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_iffalse := VAR_in28;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_iftrue := VAR_in29;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_iftrue := VAR_in3;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_iffalse := VAR_in30;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_iftrue := VAR_in31;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_iffalse := VAR_in32;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_iftrue := VAR_in33;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_iffalse := VAR_in34;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_iftrue := VAR_in35;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_iffalse := VAR_in36;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_iftrue := VAR_in37;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iffalse := VAR_in38;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iftrue := VAR_in39;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_iffalse := VAR_in4;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_iffalse := VAR_in40;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_iftrue := VAR_in41;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_iffalse := VAR_in42;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_iftrue := VAR_in43;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_iffalse := VAR_in44;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_iftrue := VAR_in45;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_iffalse := VAR_in46;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_iftrue := VAR_in47;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_iffalse := VAR_in48;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_iftrue := VAR_in49;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_iftrue := VAR_in5;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_iffalse := VAR_in50;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_iftrue := VAR_in51;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_iffalse := VAR_in52;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_iftrue := VAR_in53;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iffalse := VAR_in54;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iftrue := VAR_in55;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iffalse := VAR_in56;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iftrue := VAR_in57;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_iffalse := VAR_in58;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_iftrue := VAR_in59;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iffalse := VAR_in6;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_iffalse := VAR_in60;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_iftrue := VAR_in61;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_iffalse := VAR_in62;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_iftrue := VAR_in63;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_iffalse := VAR_in64;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_iftrue := VAR_in65;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_iffalse := VAR_in66;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_iftrue := VAR_in67;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_iffalse := VAR_in68;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_iftrue := VAR_in69;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iftrue := VAR_in7;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_iffalse := VAR_in70;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_iftrue := VAR_in71;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_iffalse := VAR_in72;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_iftrue := VAR_in73;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_iffalse := VAR_in74;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_iftrue := VAR_in75;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_iffalse := VAR_in76;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_iftrue := VAR_in77;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_iffalse := VAR_in78;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_iftrue := VAR_in79;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iffalse := VAR_in8;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_iffalse := VAR_in80;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_iftrue := VAR_in81;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_iffalse := VAR_in82;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_iftrue := VAR_in83;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_iffalse := VAR_in84;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_iftrue := VAR_in85;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_iffalse := VAR_in86;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_iftrue := VAR_in87;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_iffalse := VAR_in88;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_iftrue := VAR_in89;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iftrue := VAR_in9;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_iffalse := VAR_in90;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_iftrue := VAR_in91;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_iffalse := VAR_in92;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_iftrue := VAR_in93;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_iffalse := VAR_in94;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_iftrue := VAR_in95;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_iffalse := VAR_in96;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_iftrue := VAR_in97;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_iffalse := VAR_in98;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_iftrue := VAR_in99;
     -- uint7_2_2[bit_math_h_l1082_c10_b27d] LATENCY=0
     VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output := uint7_2_2(
     VAR_sel);

     -- uint7_0_0[bit_math_h_l14_c10_e9b9] LATENCY=0
     VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output := uint7_0_0(
     VAR_sel);

     -- uint7_6_6[bit_math_h_l1436_c10_41fb] LATENCY=0
     VAR_uint7_6_6_bit_math_h_l1436_c10_41fb_return_output := uint7_6_6(
     VAR_sel);

     -- uint7_1_1[bit_math_h_l724_c10_d539] LATENCY=0
     VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output := uint7_1_1(
     VAR_sel);

     -- uint7_3_3[bit_math_h_l1264_c10_8c95] LATENCY=0
     VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output := uint7_3_3(
     VAR_sel);

     -- uint7_4_4[bit_math_h_l1358_c10_39f5] LATENCY=0
     VAR_uint7_4_4_bit_math_h_l1358_c10_39f5_return_output := uint7_4_4(
     VAR_sel);

     -- uint7_5_5[bit_math_h_l1408_c10_5487] LATENCY=0
     VAR_uint7_5_5_bit_math_h_l1408_c10_5487_return_output := uint7_5_5(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_e9b9_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d539_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_b27d_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_8c95_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_39f5_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_39f5_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_39f5_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_39f5_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_5487_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_5487_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_cond := VAR_uint7_6_6_bit_math_h_l1436_c10_41fb_return_output;
     -- layer0_node1_MUX[bit_math_h_l29_c3_419a] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_419a_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_419a_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_419a_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output := layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output;

     -- layer0_node60_MUX[bit_math_h_l678_c3_51ce] LATENCY=0
     -- Inputs
     layer0_node60_MUX_bit_math_h_l678_c3_51ce_cond <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_cond;
     layer0_node60_MUX_bit_math_h_l678_c3_51ce_iftrue <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_iftrue;
     layer0_node60_MUX_bit_math_h_l678_c3_51ce_iffalse <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_iffalse;
     -- Outputs
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output := layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output;

     -- layer0_node33_MUX[bit_math_h_l381_c3_53ee] LATENCY=0
     -- Inputs
     layer0_node33_MUX_bit_math_h_l381_c3_53ee_cond <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_cond;
     layer0_node33_MUX_bit_math_h_l381_c3_53ee_iftrue <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_iftrue;
     layer0_node33_MUX_bit_math_h_l381_c3_53ee_iffalse <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_iffalse;
     -- Outputs
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output := layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output;

     -- layer0_node18_MUX[bit_math_h_l216_c3_6aca] LATENCY=0
     -- Inputs
     layer0_node18_MUX_bit_math_h_l216_c3_6aca_cond <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_cond;
     layer0_node18_MUX_bit_math_h_l216_c3_6aca_iftrue <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_iftrue;
     layer0_node18_MUX_bit_math_h_l216_c3_6aca_iffalse <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_iffalse;
     -- Outputs
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output := layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output;

     -- layer0_node35_MUX[bit_math_h_l403_c3_00e8] LATENCY=0
     -- Inputs
     layer0_node35_MUX_bit_math_h_l403_c3_00e8_cond <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_cond;
     layer0_node35_MUX_bit_math_h_l403_c3_00e8_iftrue <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_iftrue;
     layer0_node35_MUX_bit_math_h_l403_c3_00e8_iffalse <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_iffalse;
     -- Outputs
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output := layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output;

     -- layer0_node63_MUX[bit_math_h_l711_c3_c233] LATENCY=0
     -- Inputs
     layer0_node63_MUX_bit_math_h_l711_c3_c233_cond <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_cond;
     layer0_node63_MUX_bit_math_h_l711_c3_c233_iftrue <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_iftrue;
     layer0_node63_MUX_bit_math_h_l711_c3_c233_iffalse <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_iffalse;
     -- Outputs
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output := layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output;

     -- layer0_node17_MUX[bit_math_h_l205_c3_983c] LATENCY=0
     -- Inputs
     layer0_node17_MUX_bit_math_h_l205_c3_983c_cond <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_cond;
     layer0_node17_MUX_bit_math_h_l205_c3_983c_iftrue <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_iftrue;
     layer0_node17_MUX_bit_math_h_l205_c3_983c_iffalse <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_iffalse;
     -- Outputs
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output := layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output;

     -- layer0_node31_MUX[bit_math_h_l359_c3_a259] LATENCY=0
     -- Inputs
     layer0_node31_MUX_bit_math_h_l359_c3_a259_cond <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_cond;
     layer0_node31_MUX_bit_math_h_l359_c3_a259_iftrue <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_iftrue;
     layer0_node31_MUX_bit_math_h_l359_c3_a259_iffalse <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_iffalse;
     -- Outputs
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output := layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output;

     -- layer0_node54_MUX[bit_math_h_l612_c3_b44b] LATENCY=0
     -- Inputs
     layer0_node54_MUX_bit_math_h_l612_c3_b44b_cond <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_cond;
     layer0_node54_MUX_bit_math_h_l612_c3_b44b_iftrue <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_iftrue;
     layer0_node54_MUX_bit_math_h_l612_c3_b44b_iffalse <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_iffalse;
     -- Outputs
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output := layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output;

     -- layer0_node34_MUX[bit_math_h_l392_c3_e101] LATENCY=0
     -- Inputs
     layer0_node34_MUX_bit_math_h_l392_c3_e101_cond <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_cond;
     layer0_node34_MUX_bit_math_h_l392_c3_e101_iftrue <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_iftrue;
     layer0_node34_MUX_bit_math_h_l392_c3_e101_iffalse <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_iffalse;
     -- Outputs
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output := layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output;

     -- layer0_node9_MUX[bit_math_h_l117_c3_521d] LATENCY=0
     -- Inputs
     layer0_node9_MUX_bit_math_h_l117_c3_521d_cond <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_cond;
     layer0_node9_MUX_bit_math_h_l117_c3_521d_iftrue <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_iftrue;
     layer0_node9_MUX_bit_math_h_l117_c3_521d_iffalse <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_iffalse;
     -- Outputs
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output := layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output;

     -- layer0_node58_MUX[bit_math_h_l656_c3_485d] LATENCY=0
     -- Inputs
     layer0_node58_MUX_bit_math_h_l656_c3_485d_cond <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_cond;
     layer0_node58_MUX_bit_math_h_l656_c3_485d_iftrue <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_iftrue;
     layer0_node58_MUX_bit_math_h_l656_c3_485d_iffalse <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_iffalse;
     -- Outputs
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output := layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output;

     -- layer0_node16_MUX[bit_math_h_l194_c3_2677] LATENCY=0
     -- Inputs
     layer0_node16_MUX_bit_math_h_l194_c3_2677_cond <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_cond;
     layer0_node16_MUX_bit_math_h_l194_c3_2677_iftrue <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_iftrue;
     layer0_node16_MUX_bit_math_h_l194_c3_2677_iffalse <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_iffalse;
     -- Outputs
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output := layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output;

     -- layer0_node21_MUX[bit_math_h_l249_c3_c899] LATENCY=0
     -- Inputs
     layer0_node21_MUX_bit_math_h_l249_c3_c899_cond <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_cond;
     layer0_node21_MUX_bit_math_h_l249_c3_c899_iftrue <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_iftrue;
     layer0_node21_MUX_bit_math_h_l249_c3_c899_iffalse <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_iffalse;
     -- Outputs
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output := layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output;

     -- layer0_node10_MUX[bit_math_h_l128_c3_74ca] LATENCY=0
     -- Inputs
     layer0_node10_MUX_bit_math_h_l128_c3_74ca_cond <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_cond;
     layer0_node10_MUX_bit_math_h_l128_c3_74ca_iftrue <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_iftrue;
     layer0_node10_MUX_bit_math_h_l128_c3_74ca_iffalse <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_iffalse;
     -- Outputs
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output := layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output;

     -- layer0_node40_MUX[bit_math_h_l458_c3_0262] LATENCY=0
     -- Inputs
     layer0_node40_MUX_bit_math_h_l458_c3_0262_cond <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_cond;
     layer0_node40_MUX_bit_math_h_l458_c3_0262_iftrue <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_iftrue;
     layer0_node40_MUX_bit_math_h_l458_c3_0262_iffalse <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_iffalse;
     -- Outputs
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output := layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output;

     -- layer0_node12_MUX[bit_math_h_l150_c3_ce47] LATENCY=0
     -- Inputs
     layer0_node12_MUX_bit_math_h_l150_c3_ce47_cond <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_cond;
     layer0_node12_MUX_bit_math_h_l150_c3_ce47_iftrue <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_iftrue;
     layer0_node12_MUX_bit_math_h_l150_c3_ce47_iffalse <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_iffalse;
     -- Outputs
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output := layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output;

     -- layer0_node20_MUX[bit_math_h_l238_c3_27b2] LATENCY=0
     -- Inputs
     layer0_node20_MUX_bit_math_h_l238_c3_27b2_cond <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_cond;
     layer0_node20_MUX_bit_math_h_l238_c3_27b2_iftrue <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_iftrue;
     layer0_node20_MUX_bit_math_h_l238_c3_27b2_iffalse <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_iffalse;
     -- Outputs
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output := layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output;

     -- layer0_node49_MUX[bit_math_h_l557_c3_44e2] LATENCY=0
     -- Inputs
     layer0_node49_MUX_bit_math_h_l557_c3_44e2_cond <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_cond;
     layer0_node49_MUX_bit_math_h_l557_c3_44e2_iftrue <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_iftrue;
     layer0_node49_MUX_bit_math_h_l557_c3_44e2_iffalse <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_iffalse;
     -- Outputs
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output := layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output;

     -- layer0_node56_MUX[bit_math_h_l634_c3_6313] LATENCY=0
     -- Inputs
     layer0_node56_MUX_bit_math_h_l634_c3_6313_cond <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_cond;
     layer0_node56_MUX_bit_math_h_l634_c3_6313_iftrue <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_iftrue;
     layer0_node56_MUX_bit_math_h_l634_c3_6313_iffalse <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_iffalse;
     -- Outputs
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output := layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_7a6b] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_7a6b_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output := layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output;

     -- layer0_node8_MUX[bit_math_h_l106_c3_0c54] LATENCY=0
     -- Inputs
     layer0_node8_MUX_bit_math_h_l106_c3_0c54_cond <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_cond;
     layer0_node8_MUX_bit_math_h_l106_c3_0c54_iftrue <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_iftrue;
     layer0_node8_MUX_bit_math_h_l106_c3_0c54_iffalse <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_iffalse;
     -- Outputs
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output := layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_1ccf] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_1ccf_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output := layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output;

     -- layer0_node57_MUX[bit_math_h_l645_c3_d8b1] LATENCY=0
     -- Inputs
     layer0_node57_MUX_bit_math_h_l645_c3_d8b1_cond <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_cond;
     layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iftrue <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iftrue;
     layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iffalse <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_iffalse;
     -- Outputs
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output := layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output;

     -- layer0_node15_MUX[bit_math_h_l183_c3_d015] LATENCY=0
     -- Inputs
     layer0_node15_MUX_bit_math_h_l183_c3_d015_cond <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_cond;
     layer0_node15_MUX_bit_math_h_l183_c3_d015_iftrue <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_iftrue;
     layer0_node15_MUX_bit_math_h_l183_c3_d015_iffalse <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_iffalse;
     -- Outputs
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output := layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output;

     -- layer0_node36_MUX[bit_math_h_l414_c3_d477] LATENCY=0
     -- Inputs
     layer0_node36_MUX_bit_math_h_l414_c3_d477_cond <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_cond;
     layer0_node36_MUX_bit_math_h_l414_c3_d477_iftrue <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_iftrue;
     layer0_node36_MUX_bit_math_h_l414_c3_d477_iffalse <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_iffalse;
     -- Outputs
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output := layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output;

     -- layer0_node46_MUX[bit_math_h_l524_c3_1b28] LATENCY=0
     -- Inputs
     layer0_node46_MUX_bit_math_h_l524_c3_1b28_cond <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_cond;
     layer0_node46_MUX_bit_math_h_l524_c3_1b28_iftrue <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_iftrue;
     layer0_node46_MUX_bit_math_h_l524_c3_1b28_iffalse <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_iffalse;
     -- Outputs
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output := layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_ffca] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_ffca_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_ffca_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_ffca_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output := layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output;

     -- layer0_node47_MUX[bit_math_h_l535_c3_8ede] LATENCY=0
     -- Inputs
     layer0_node47_MUX_bit_math_h_l535_c3_8ede_cond <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_cond;
     layer0_node47_MUX_bit_math_h_l535_c3_8ede_iftrue <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_iftrue;
     layer0_node47_MUX_bit_math_h_l535_c3_8ede_iffalse <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_iffalse;
     -- Outputs
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output := layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output;

     -- layer0_node42_MUX[bit_math_h_l480_c3_45fb] LATENCY=0
     -- Inputs
     layer0_node42_MUX_bit_math_h_l480_c3_45fb_cond <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_cond;
     layer0_node42_MUX_bit_math_h_l480_c3_45fb_iftrue <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_iftrue;
     layer0_node42_MUX_bit_math_h_l480_c3_45fb_iffalse <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_iffalse;
     -- Outputs
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output := layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output;

     -- layer0_node22_MUX[bit_math_h_l260_c3_0382] LATENCY=0
     -- Inputs
     layer0_node22_MUX_bit_math_h_l260_c3_0382_cond <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_cond;
     layer0_node22_MUX_bit_math_h_l260_c3_0382_iftrue <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_iftrue;
     layer0_node22_MUX_bit_math_h_l260_c3_0382_iffalse <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_iffalse;
     -- Outputs
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output := layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output;

     -- layer0_node51_MUX[bit_math_h_l579_c3_a08f] LATENCY=0
     -- Inputs
     layer0_node51_MUX_bit_math_h_l579_c3_a08f_cond <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_cond;
     layer0_node51_MUX_bit_math_h_l579_c3_a08f_iftrue <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_iftrue;
     layer0_node51_MUX_bit_math_h_l579_c3_a08f_iffalse <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_iffalse;
     -- Outputs
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output := layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output;

     -- layer0_node30_MUX[bit_math_h_l348_c3_c538] LATENCY=0
     -- Inputs
     layer0_node30_MUX_bit_math_h_l348_c3_c538_cond <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_cond;
     layer0_node30_MUX_bit_math_h_l348_c3_c538_iftrue <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_iftrue;
     layer0_node30_MUX_bit_math_h_l348_c3_c538_iffalse <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_iffalse;
     -- Outputs
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output := layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output;

     -- layer0_node52_MUX[bit_math_h_l590_c3_f2e8] LATENCY=0
     -- Inputs
     layer0_node52_MUX_bit_math_h_l590_c3_f2e8_cond <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_cond;
     layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iftrue <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iftrue;
     layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iffalse <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_iffalse;
     -- Outputs
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output := layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output;

     -- layer0_node26_MUX[bit_math_h_l304_c3_53c3] LATENCY=0
     -- Inputs
     layer0_node26_MUX_bit_math_h_l304_c3_53c3_cond <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_cond;
     layer0_node26_MUX_bit_math_h_l304_c3_53c3_iftrue <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_iftrue;
     layer0_node26_MUX_bit_math_h_l304_c3_53c3_iffalse <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_iffalse;
     -- Outputs
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output := layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output;

     -- layer0_node61_MUX[bit_math_h_l689_c3_8d98] LATENCY=0
     -- Inputs
     layer0_node61_MUX_bit_math_h_l689_c3_8d98_cond <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_cond;
     layer0_node61_MUX_bit_math_h_l689_c3_8d98_iftrue <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_iftrue;
     layer0_node61_MUX_bit_math_h_l689_c3_8d98_iffalse <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_iffalse;
     -- Outputs
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output := layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_5094] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_5094_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_5094_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_5094_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output := layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_0dd3] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_0dd3_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output := layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output;

     -- layer0_node45_MUX[bit_math_h_l513_c3_405f] LATENCY=0
     -- Inputs
     layer0_node45_MUX_bit_math_h_l513_c3_405f_cond <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_cond;
     layer0_node45_MUX_bit_math_h_l513_c3_405f_iftrue <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_iftrue;
     layer0_node45_MUX_bit_math_h_l513_c3_405f_iffalse <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_iffalse;
     -- Outputs
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output := layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output;

     -- layer0_node24_MUX[bit_math_h_l282_c3_de03] LATENCY=0
     -- Inputs
     layer0_node24_MUX_bit_math_h_l282_c3_de03_cond <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_cond;
     layer0_node24_MUX_bit_math_h_l282_c3_de03_iftrue <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_iftrue;
     layer0_node24_MUX_bit_math_h_l282_c3_de03_iffalse <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_iffalse;
     -- Outputs
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output := layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output;

     -- layer0_node28_MUX[bit_math_h_l326_c3_a3f6] LATENCY=0
     -- Inputs
     layer0_node28_MUX_bit_math_h_l326_c3_a3f6_cond <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_cond;
     layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iftrue <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iftrue;
     layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iffalse <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_iffalse;
     -- Outputs
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output := layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output;

     -- layer0_node53_MUX[bit_math_h_l601_c3_33d0] LATENCY=0
     -- Inputs
     layer0_node53_MUX_bit_math_h_l601_c3_33d0_cond <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_cond;
     layer0_node53_MUX_bit_math_h_l601_c3_33d0_iftrue <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_iftrue;
     layer0_node53_MUX_bit_math_h_l601_c3_33d0_iffalse <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_iffalse;
     -- Outputs
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output := layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output;

     -- layer0_node55_MUX[bit_math_h_l623_c3_0aaf] LATENCY=0
     -- Inputs
     layer0_node55_MUX_bit_math_h_l623_c3_0aaf_cond <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_cond;
     layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iftrue <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iftrue;
     layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iffalse <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_iffalse;
     -- Outputs
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output := layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output;

     -- layer0_node43_MUX[bit_math_h_l491_c3_0137] LATENCY=0
     -- Inputs
     layer0_node43_MUX_bit_math_h_l491_c3_0137_cond <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_cond;
     layer0_node43_MUX_bit_math_h_l491_c3_0137_iftrue <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_iftrue;
     layer0_node43_MUX_bit_math_h_l491_c3_0137_iffalse <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_iffalse;
     -- Outputs
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output := layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output;

     -- layer0_node39_MUX[bit_math_h_l447_c3_50eb] LATENCY=0
     -- Inputs
     layer0_node39_MUX_bit_math_h_l447_c3_50eb_cond <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_cond;
     layer0_node39_MUX_bit_math_h_l447_c3_50eb_iftrue <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_iftrue;
     layer0_node39_MUX_bit_math_h_l447_c3_50eb_iffalse <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_iffalse;
     -- Outputs
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output := layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output;

     -- layer0_node25_MUX[bit_math_h_l293_c3_32f2] LATENCY=0
     -- Inputs
     layer0_node25_MUX_bit_math_h_l293_c3_32f2_cond <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_cond;
     layer0_node25_MUX_bit_math_h_l293_c3_32f2_iftrue <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_iftrue;
     layer0_node25_MUX_bit_math_h_l293_c3_32f2_iffalse <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_iffalse;
     -- Outputs
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output := layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output;

     -- layer0_node44_MUX[bit_math_h_l502_c3_983c] LATENCY=0
     -- Inputs
     layer0_node44_MUX_bit_math_h_l502_c3_983c_cond <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_cond;
     layer0_node44_MUX_bit_math_h_l502_c3_983c_iftrue <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_iftrue;
     layer0_node44_MUX_bit_math_h_l502_c3_983c_iffalse <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_iffalse;
     -- Outputs
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output := layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output;

     -- layer0_node19_MUX[bit_math_h_l227_c3_1ba6] LATENCY=0
     -- Inputs
     layer0_node19_MUX_bit_math_h_l227_c3_1ba6_cond <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_cond;
     layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iftrue <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iftrue;
     layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iffalse <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_iffalse;
     -- Outputs
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output := layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output;

     -- layer0_node38_MUX[bit_math_h_l436_c3_0345] LATENCY=0
     -- Inputs
     layer0_node38_MUX_bit_math_h_l436_c3_0345_cond <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_cond;
     layer0_node38_MUX_bit_math_h_l436_c3_0345_iftrue <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_iftrue;
     layer0_node38_MUX_bit_math_h_l436_c3_0345_iffalse <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_iffalse;
     -- Outputs
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output := layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output;

     -- layer0_node41_MUX[bit_math_h_l469_c3_4656] LATENCY=0
     -- Inputs
     layer0_node41_MUX_bit_math_h_l469_c3_4656_cond <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_cond;
     layer0_node41_MUX_bit_math_h_l469_c3_4656_iftrue <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_iftrue;
     layer0_node41_MUX_bit_math_h_l469_c3_4656_iffalse <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_iffalse;
     -- Outputs
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output := layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output;

     -- layer0_node59_MUX[bit_math_h_l667_c3_6892] LATENCY=0
     -- Inputs
     layer0_node59_MUX_bit_math_h_l667_c3_6892_cond <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_cond;
     layer0_node59_MUX_bit_math_h_l667_c3_6892_iftrue <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_iftrue;
     layer0_node59_MUX_bit_math_h_l667_c3_6892_iffalse <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_iffalse;
     -- Outputs
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output := layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output;

     -- layer0_node23_MUX[bit_math_h_l271_c3_93d7] LATENCY=0
     -- Inputs
     layer0_node23_MUX_bit_math_h_l271_c3_93d7_cond <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_cond;
     layer0_node23_MUX_bit_math_h_l271_c3_93d7_iftrue <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_iftrue;
     layer0_node23_MUX_bit_math_h_l271_c3_93d7_iffalse <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_iffalse;
     -- Outputs
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output := layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output;

     -- layer0_node13_MUX[bit_math_h_l161_c3_76bd] LATENCY=0
     -- Inputs
     layer0_node13_MUX_bit_math_h_l161_c3_76bd_cond <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_cond;
     layer0_node13_MUX_bit_math_h_l161_c3_76bd_iftrue <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_iftrue;
     layer0_node13_MUX_bit_math_h_l161_c3_76bd_iffalse <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_iffalse;
     -- Outputs
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output := layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output;

     -- layer0_node11_MUX[bit_math_h_l139_c3_31b7] LATENCY=0
     -- Inputs
     layer0_node11_MUX_bit_math_h_l139_c3_31b7_cond <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_cond;
     layer0_node11_MUX_bit_math_h_l139_c3_31b7_iftrue <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_iftrue;
     layer0_node11_MUX_bit_math_h_l139_c3_31b7_iffalse <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_iffalse;
     -- Outputs
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output := layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_195c] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_195c_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_195c_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_195c_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output := layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output;

     -- layer0_node14_MUX[bit_math_h_l172_c3_7b21] LATENCY=0
     -- Inputs
     layer0_node14_MUX_bit_math_h_l172_c3_7b21_cond <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_cond;
     layer0_node14_MUX_bit_math_h_l172_c3_7b21_iftrue <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_iftrue;
     layer0_node14_MUX_bit_math_h_l172_c3_7b21_iffalse <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_iffalse;
     -- Outputs
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output := layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output;

     -- layer0_node29_MUX[bit_math_h_l337_c3_76ce] LATENCY=0
     -- Inputs
     layer0_node29_MUX_bit_math_h_l337_c3_76ce_cond <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_cond;
     layer0_node29_MUX_bit_math_h_l337_c3_76ce_iftrue <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_iftrue;
     layer0_node29_MUX_bit_math_h_l337_c3_76ce_iffalse <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_iffalse;
     -- Outputs
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output := layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output;

     -- layer0_node48_MUX[bit_math_h_l546_c3_f942] LATENCY=0
     -- Inputs
     layer0_node48_MUX_bit_math_h_l546_c3_f942_cond <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_cond;
     layer0_node48_MUX_bit_math_h_l546_c3_f942_iftrue <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_iftrue;
     layer0_node48_MUX_bit_math_h_l546_c3_f942_iffalse <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_iffalse;
     -- Outputs
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output := layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output;

     -- layer0_node50_MUX[bit_math_h_l568_c3_1207] LATENCY=0
     -- Inputs
     layer0_node50_MUX_bit_math_h_l568_c3_1207_cond <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_cond;
     layer0_node50_MUX_bit_math_h_l568_c3_1207_iftrue <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_iftrue;
     layer0_node50_MUX_bit_math_h_l568_c3_1207_iffalse <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_iffalse;
     -- Outputs
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output := layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output;

     -- layer0_node37_MUX[bit_math_h_l425_c3_bb07] LATENCY=0
     -- Inputs
     layer0_node37_MUX_bit_math_h_l425_c3_bb07_cond <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_cond;
     layer0_node37_MUX_bit_math_h_l425_c3_bb07_iftrue <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_iftrue;
     layer0_node37_MUX_bit_math_h_l425_c3_bb07_iffalse <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_iffalse;
     -- Outputs
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output := layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output;

     -- layer0_node62_MUX[bit_math_h_l700_c3_9327] LATENCY=0
     -- Inputs
     layer0_node62_MUX_bit_math_h_l700_c3_9327_cond <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_cond;
     layer0_node62_MUX_bit_math_h_l700_c3_9327_iftrue <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_iftrue;
     layer0_node62_MUX_bit_math_h_l700_c3_9327_iffalse <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_iffalse;
     -- Outputs
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output := layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output;

     -- layer0_node27_MUX[bit_math_h_l315_c3_e4a1] LATENCY=0
     -- Inputs
     layer0_node27_MUX_bit_math_h_l315_c3_e4a1_cond <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_cond;
     layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iftrue <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iftrue;
     layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iffalse <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_iffalse;
     -- Outputs
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output := layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output;

     -- layer0_node32_MUX[bit_math_h_l370_c3_2900] LATENCY=0
     -- Inputs
     layer0_node32_MUX_bit_math_h_l370_c3_2900_cond <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_cond;
     layer0_node32_MUX_bit_math_h_l370_c3_2900_iftrue <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_iftrue;
     layer0_node32_MUX_bit_math_h_l370_c3_2900_iffalse <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_iffalse;
     -- Outputs
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output := layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_7e59] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_7e59_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_7e59_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_7e59_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output := layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_5094_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_iffalse := VAR_layer0_node10_MUX_bit_math_h_l128_c3_74ca_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_iftrue := VAR_layer0_node11_MUX_bit_math_h_l139_c3_31b7_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_iffalse := VAR_layer0_node12_MUX_bit_math_h_l150_c3_ce47_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_iftrue := VAR_layer0_node13_MUX_bit_math_h_l161_c3_76bd_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_iffalse := VAR_layer0_node14_MUX_bit_math_h_l172_c3_7b21_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_iftrue := VAR_layer0_node15_MUX_bit_math_h_l183_c3_d015_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_iffalse := VAR_layer0_node16_MUX_bit_math_h_l194_c3_2677_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_iftrue := VAR_layer0_node17_MUX_bit_math_h_l205_c3_983c_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iffalse := VAR_layer0_node18_MUX_bit_math_h_l216_c3_6aca_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iftrue := VAR_layer0_node19_MUX_bit_math_h_l227_c3_1ba6_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_419a_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iffalse := VAR_layer0_node20_MUX_bit_math_h_l238_c3_27b2_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iftrue := VAR_layer0_node21_MUX_bit_math_h_l249_c3_c899_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iffalse := VAR_layer0_node22_MUX_bit_math_h_l260_c3_0382_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iftrue := VAR_layer0_node23_MUX_bit_math_h_l271_c3_93d7_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_iffalse := VAR_layer0_node24_MUX_bit_math_h_l282_c3_de03_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_iftrue := VAR_layer0_node25_MUX_bit_math_h_l293_c3_32f2_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_iffalse := VAR_layer0_node26_MUX_bit_math_h_l304_c3_53c3_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_iftrue := VAR_layer0_node27_MUX_bit_math_h_l315_c3_e4a1_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_iffalse := VAR_layer0_node28_MUX_bit_math_h_l326_c3_a3f6_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_iftrue := VAR_layer0_node29_MUX_bit_math_h_l337_c3_76ce_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_195c_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iffalse := VAR_layer0_node30_MUX_bit_math_h_l348_c3_c538_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iftrue := VAR_layer0_node31_MUX_bit_math_h_l359_c3_a259_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_iffalse := VAR_layer0_node32_MUX_bit_math_h_l370_c3_2900_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_iftrue := VAR_layer0_node33_MUX_bit_math_h_l381_c3_53ee_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_iffalse := VAR_layer0_node34_MUX_bit_math_h_l392_c3_e101_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_iftrue := VAR_layer0_node35_MUX_bit_math_h_l403_c3_00e8_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iffalse := VAR_layer0_node36_MUX_bit_math_h_l414_c3_d477_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iftrue := VAR_layer0_node37_MUX_bit_math_h_l425_c3_bb07_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_iffalse := VAR_layer0_node38_MUX_bit_math_h_l436_c3_0345_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_iftrue := VAR_layer0_node39_MUX_bit_math_h_l447_c3_50eb_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_7a6b_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_iffalse := VAR_layer0_node40_MUX_bit_math_h_l458_c3_0262_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_iftrue := VAR_layer0_node41_MUX_bit_math_h_l469_c3_4656_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_iffalse := VAR_layer0_node42_MUX_bit_math_h_l480_c3_45fb_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_iftrue := VAR_layer0_node43_MUX_bit_math_h_l491_c3_0137_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_iffalse := VAR_layer0_node44_MUX_bit_math_h_l502_c3_983c_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_iftrue := VAR_layer0_node45_MUX_bit_math_h_l513_c3_405f_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_iffalse := VAR_layer0_node46_MUX_bit_math_h_l524_c3_1b28_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_iftrue := VAR_layer0_node47_MUX_bit_math_h_l535_c3_8ede_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iffalse := VAR_layer0_node48_MUX_bit_math_h_l546_c3_f942_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iftrue := VAR_layer0_node49_MUX_bit_math_h_l557_c3_44e2_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_1ccf_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_iffalse := VAR_layer0_node50_MUX_bit_math_h_l568_c3_1207_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_iftrue := VAR_layer0_node51_MUX_bit_math_h_l579_c3_a08f_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iffalse := VAR_layer0_node52_MUX_bit_math_h_l590_c3_f2e8_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iftrue := VAR_layer0_node53_MUX_bit_math_h_l601_c3_33d0_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iffalse := VAR_layer0_node54_MUX_bit_math_h_l612_c3_b44b_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iftrue := VAR_layer0_node55_MUX_bit_math_h_l623_c3_0aaf_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_iffalse := VAR_layer0_node56_MUX_bit_math_h_l634_c3_6313_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_iftrue := VAR_layer0_node57_MUX_bit_math_h_l645_c3_d8b1_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_iffalse := VAR_layer0_node58_MUX_bit_math_h_l656_c3_485d_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_iftrue := VAR_layer0_node59_MUX_bit_math_h_l667_c3_6892_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_0dd3_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iffalse := VAR_layer0_node60_MUX_bit_math_h_l678_c3_51ce_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iftrue := VAR_layer0_node61_MUX_bit_math_h_l689_c3_8d98_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_iffalse := VAR_layer0_node62_MUX_bit_math_h_l700_c3_9327_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_iftrue := VAR_layer0_node63_MUX_bit_math_h_l711_c3_c233_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_7e59_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_ffca_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_iffalse := VAR_layer0_node8_MUX_bit_math_h_l106_c3_0c54_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_iftrue := VAR_layer0_node9_MUX_bit_math_h_l117_c3_521d_return_output;
     -- layer1_node22_MUX[bit_math_h_l970_c3_8998] LATENCY=0
     -- Inputs
     layer1_node22_MUX_bit_math_h_l970_c3_8998_cond <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_cond;
     layer1_node22_MUX_bit_math_h_l970_c3_8998_iftrue <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_iftrue;
     layer1_node22_MUX_bit_math_h_l970_c3_8998_iffalse <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_iffalse;
     -- Outputs
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output := layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output;

     -- layer1_node20_MUX[bit_math_h_l948_c3_2d00] LATENCY=0
     -- Inputs
     layer1_node20_MUX_bit_math_h_l948_c3_2d00_cond <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_cond;
     layer1_node20_MUX_bit_math_h_l948_c3_2d00_iftrue <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_iftrue;
     layer1_node20_MUX_bit_math_h_l948_c3_2d00_iffalse <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_iffalse;
     -- Outputs
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output := layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output;

     -- layer1_node31_MUX[bit_math_h_l1069_c3_5488] LATENCY=0
     -- Inputs
     layer1_node31_MUX_bit_math_h_l1069_c3_5488_cond <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_cond;
     layer1_node31_MUX_bit_math_h_l1069_c3_5488_iftrue <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_iftrue;
     layer1_node31_MUX_bit_math_h_l1069_c3_5488_iffalse <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_iffalse;
     -- Outputs
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output := layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output;

     -- layer1_node4_MUX[bit_math_h_l772_c3_a071] LATENCY=0
     -- Inputs
     layer1_node4_MUX_bit_math_h_l772_c3_a071_cond <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_cond;
     layer1_node4_MUX_bit_math_h_l772_c3_a071_iftrue <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_iftrue;
     layer1_node4_MUX_bit_math_h_l772_c3_a071_iffalse <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_iffalse;
     -- Outputs
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output := layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output;

     -- layer1_node11_MUX[bit_math_h_l849_c3_2cb0] LATENCY=0
     -- Inputs
     layer1_node11_MUX_bit_math_h_l849_c3_2cb0_cond <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_cond;
     layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iftrue <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iftrue;
     layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iffalse <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_iffalse;
     -- Outputs
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output := layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output;

     -- layer1_node17_MUX[bit_math_h_l915_c3_90a2] LATENCY=0
     -- Inputs
     layer1_node17_MUX_bit_math_h_l915_c3_90a2_cond <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_cond;
     layer1_node17_MUX_bit_math_h_l915_c3_90a2_iftrue <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_iftrue;
     layer1_node17_MUX_bit_math_h_l915_c3_90a2_iffalse <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_iffalse;
     -- Outputs
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output := layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output;

     -- layer1_node26_MUX[bit_math_h_l1014_c3_1e7d] LATENCY=0
     -- Inputs
     layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_cond <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_cond;
     layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iftrue <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iftrue;
     layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iffalse <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_iffalse;
     -- Outputs
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output := layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output;

     -- layer1_node23_MUX[bit_math_h_l981_c3_102a] LATENCY=0
     -- Inputs
     layer1_node23_MUX_bit_math_h_l981_c3_102a_cond <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_cond;
     layer1_node23_MUX_bit_math_h_l981_c3_102a_iftrue <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_iftrue;
     layer1_node23_MUX_bit_math_h_l981_c3_102a_iffalse <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_iffalse;
     -- Outputs
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output := layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output;

     -- layer1_node8_MUX[bit_math_h_l816_c3_fa37] LATENCY=0
     -- Inputs
     layer1_node8_MUX_bit_math_h_l816_c3_fa37_cond <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_cond;
     layer1_node8_MUX_bit_math_h_l816_c3_fa37_iftrue <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_iftrue;
     layer1_node8_MUX_bit_math_h_l816_c3_fa37_iffalse <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_iffalse;
     -- Outputs
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output := layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output;

     -- layer1_node16_MUX[bit_math_h_l904_c3_234e] LATENCY=0
     -- Inputs
     layer1_node16_MUX_bit_math_h_l904_c3_234e_cond <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_cond;
     layer1_node16_MUX_bit_math_h_l904_c3_234e_iftrue <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_iftrue;
     layer1_node16_MUX_bit_math_h_l904_c3_234e_iffalse <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_iffalse;
     -- Outputs
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output := layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output;

     -- layer1_node29_MUX[bit_math_h_l1047_c3_3314] LATENCY=0
     -- Inputs
     layer1_node29_MUX_bit_math_h_l1047_c3_3314_cond <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_cond;
     layer1_node29_MUX_bit_math_h_l1047_c3_3314_iftrue <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_iftrue;
     layer1_node29_MUX_bit_math_h_l1047_c3_3314_iffalse <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_iffalse;
     -- Outputs
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output := layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output;

     -- layer1_node30_MUX[bit_math_h_l1058_c3_6a5f] LATENCY=0
     -- Inputs
     layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_cond <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_cond;
     layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iftrue <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iftrue;
     layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iffalse <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_iffalse;
     -- Outputs
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output := layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output;

     -- layer1_node1_MUX[bit_math_h_l739_c3_e269] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l739_c3_e269_cond <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_cond;
     layer1_node1_MUX_bit_math_h_l739_c3_e269_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_iftrue;
     layer1_node1_MUX_bit_math_h_l739_c3_e269_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output := layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output;

     -- layer1_node15_MUX[bit_math_h_l893_c3_5e2b] LATENCY=0
     -- Inputs
     layer1_node15_MUX_bit_math_h_l893_c3_5e2b_cond <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_cond;
     layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iftrue <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iftrue;
     layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iffalse <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_iffalse;
     -- Outputs
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output := layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output;

     -- layer1_node14_MUX[bit_math_h_l882_c3_3e12] LATENCY=0
     -- Inputs
     layer1_node14_MUX_bit_math_h_l882_c3_3e12_cond <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_cond;
     layer1_node14_MUX_bit_math_h_l882_c3_3e12_iftrue <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_iftrue;
     layer1_node14_MUX_bit_math_h_l882_c3_3e12_iffalse <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_iffalse;
     -- Outputs
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output := layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output;

     -- layer1_node10_MUX[bit_math_h_l838_c3_7eb8] LATENCY=0
     -- Inputs
     layer1_node10_MUX_bit_math_h_l838_c3_7eb8_cond <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_cond;
     layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iftrue <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iftrue;
     layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iffalse <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_iffalse;
     -- Outputs
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output := layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output;

     -- layer1_node7_MUX[bit_math_h_l805_c3_c99c] LATENCY=0
     -- Inputs
     layer1_node7_MUX_bit_math_h_l805_c3_c99c_cond <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_cond;
     layer1_node7_MUX_bit_math_h_l805_c3_c99c_iftrue <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_iftrue;
     layer1_node7_MUX_bit_math_h_l805_c3_c99c_iffalse <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_iffalse;
     -- Outputs
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output := layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output;

     -- layer1_node21_MUX[bit_math_h_l959_c3_f682] LATENCY=0
     -- Inputs
     layer1_node21_MUX_bit_math_h_l959_c3_f682_cond <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_cond;
     layer1_node21_MUX_bit_math_h_l959_c3_f682_iftrue <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_iftrue;
     layer1_node21_MUX_bit_math_h_l959_c3_f682_iffalse <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_iffalse;
     -- Outputs
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output := layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output;

     -- layer1_node5_MUX[bit_math_h_l783_c3_9883] LATENCY=0
     -- Inputs
     layer1_node5_MUX_bit_math_h_l783_c3_9883_cond <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_cond;
     layer1_node5_MUX_bit_math_h_l783_c3_9883_iftrue <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_iftrue;
     layer1_node5_MUX_bit_math_h_l783_c3_9883_iffalse <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_iffalse;
     -- Outputs
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output := layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output;

     -- layer1_node2_MUX[bit_math_h_l750_c3_5aa6] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l750_c3_5aa6_cond <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_cond;
     layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iftrue;
     layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output := layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output;

     -- layer1_node18_MUX[bit_math_h_l926_c3_ecc8] LATENCY=0
     -- Inputs
     layer1_node18_MUX_bit_math_h_l926_c3_ecc8_cond <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_cond;
     layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iftrue <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iftrue;
     layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iffalse <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_iffalse;
     -- Outputs
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output := layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output;

     -- layer1_node24_MUX[bit_math_h_l992_c3_9fd6] LATENCY=0
     -- Inputs
     layer1_node24_MUX_bit_math_h_l992_c3_9fd6_cond <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_cond;
     layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iftrue <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iftrue;
     layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iffalse <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_iffalse;
     -- Outputs
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output := layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output;

     -- layer1_node9_MUX[bit_math_h_l827_c3_d6c2] LATENCY=0
     -- Inputs
     layer1_node9_MUX_bit_math_h_l827_c3_d6c2_cond <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_cond;
     layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iftrue <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iftrue;
     layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iffalse <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_iffalse;
     -- Outputs
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output := layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output;

     -- layer1_node6_MUX[bit_math_h_l794_c3_cf43] LATENCY=0
     -- Inputs
     layer1_node6_MUX_bit_math_h_l794_c3_cf43_cond <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_cond;
     layer1_node6_MUX_bit_math_h_l794_c3_cf43_iftrue <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_iftrue;
     layer1_node6_MUX_bit_math_h_l794_c3_cf43_iffalse <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_iffalse;
     -- Outputs
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output := layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output;

     -- layer1_node27_MUX[bit_math_h_l1025_c3_46dd] LATENCY=0
     -- Inputs
     layer1_node27_MUX_bit_math_h_l1025_c3_46dd_cond <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_cond;
     layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iftrue <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iftrue;
     layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iffalse <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_iffalse;
     -- Outputs
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output := layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output;

     -- layer1_node19_MUX[bit_math_h_l937_c3_7211] LATENCY=0
     -- Inputs
     layer1_node19_MUX_bit_math_h_l937_c3_7211_cond <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_cond;
     layer1_node19_MUX_bit_math_h_l937_c3_7211_iftrue <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_iftrue;
     layer1_node19_MUX_bit_math_h_l937_c3_7211_iffalse <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_iffalse;
     -- Outputs
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output := layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output;

     -- layer1_node12_MUX[bit_math_h_l860_c3_32ef] LATENCY=0
     -- Inputs
     layer1_node12_MUX_bit_math_h_l860_c3_32ef_cond <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_cond;
     layer1_node12_MUX_bit_math_h_l860_c3_32ef_iftrue <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_iftrue;
     layer1_node12_MUX_bit_math_h_l860_c3_32ef_iffalse <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_iffalse;
     -- Outputs
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output := layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output;

     -- layer1_node13_MUX[bit_math_h_l871_c3_c37d] LATENCY=0
     -- Inputs
     layer1_node13_MUX_bit_math_h_l871_c3_c37d_cond <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_cond;
     layer1_node13_MUX_bit_math_h_l871_c3_c37d_iftrue <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_iftrue;
     layer1_node13_MUX_bit_math_h_l871_c3_c37d_iffalse <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_iffalse;
     -- Outputs
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output := layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output;

     -- layer1_node28_MUX[bit_math_h_l1036_c3_4035] LATENCY=0
     -- Inputs
     layer1_node28_MUX_bit_math_h_l1036_c3_4035_cond <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_cond;
     layer1_node28_MUX_bit_math_h_l1036_c3_4035_iftrue <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_iftrue;
     layer1_node28_MUX_bit_math_h_l1036_c3_4035_iffalse <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_iffalse;
     -- Outputs
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output := layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output;

     -- layer1_node3_MUX[bit_math_h_l761_c3_850a] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l761_c3_850a_cond <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_cond;
     layer1_node3_MUX_bit_math_h_l761_c3_850a_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_iftrue;
     layer1_node3_MUX_bit_math_h_l761_c3_850a_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output := layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output;

     -- layer1_node25_MUX[bit_math_h_l1003_c3_271e] LATENCY=0
     -- Inputs
     layer1_node25_MUX_bit_math_h_l1003_c3_271e_cond <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_cond;
     layer1_node25_MUX_bit_math_h_l1003_c3_271e_iftrue <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_iftrue;
     layer1_node25_MUX_bit_math_h_l1003_c3_271e_iffalse <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_iffalse;
     -- Outputs
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output := layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output;

     -- layer1_node0_MUX[bit_math_h_l728_c3_cd45] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l728_c3_cd45_cond <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_cond;
     layer1_node0_MUX_bit_math_h_l728_c3_cd45_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_iftrue;
     layer1_node0_MUX_bit_math_h_l728_c3_cd45_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output := layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_iffalse := VAR_layer1_node0_MUX_bit_math_h_l728_c3_cd45_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iffalse := VAR_layer1_node10_MUX_bit_math_h_l838_c3_7eb8_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iftrue := VAR_layer1_node11_MUX_bit_math_h_l849_c3_2cb0_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_iffalse := VAR_layer1_node12_MUX_bit_math_h_l860_c3_32ef_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_iftrue := VAR_layer1_node13_MUX_bit_math_h_l871_c3_c37d_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iffalse := VAR_layer1_node14_MUX_bit_math_h_l882_c3_3e12_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iftrue := VAR_layer1_node15_MUX_bit_math_h_l893_c3_5e2b_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iffalse := VAR_layer1_node16_MUX_bit_math_h_l904_c3_234e_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iftrue := VAR_layer1_node17_MUX_bit_math_h_l915_c3_90a2_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iffalse := VAR_layer1_node18_MUX_bit_math_h_l926_c3_ecc8_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iftrue := VAR_layer1_node19_MUX_bit_math_h_l937_c3_7211_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_iftrue := VAR_layer1_node1_MUX_bit_math_h_l739_c3_e269_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_iffalse := VAR_layer1_node20_MUX_bit_math_h_l948_c3_2d00_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_iftrue := VAR_layer1_node21_MUX_bit_math_h_l959_c3_f682_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iffalse := VAR_layer1_node22_MUX_bit_math_h_l970_c3_8998_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iftrue := VAR_layer1_node23_MUX_bit_math_h_l981_c3_102a_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iffalse := VAR_layer1_node24_MUX_bit_math_h_l992_c3_9fd6_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iftrue := VAR_layer1_node25_MUX_bit_math_h_l1003_c3_271e_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_iffalse := VAR_layer1_node26_MUX_bit_math_h_l1014_c3_1e7d_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_iftrue := VAR_layer1_node27_MUX_bit_math_h_l1025_c3_46dd_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_iffalse := VAR_layer1_node28_MUX_bit_math_h_l1036_c3_4035_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_iftrue := VAR_layer1_node29_MUX_bit_math_h_l1047_c3_3314_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_iffalse := VAR_layer1_node2_MUX_bit_math_h_l750_c3_5aa6_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_iffalse := VAR_layer1_node30_MUX_bit_math_h_l1058_c3_6a5f_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_iftrue := VAR_layer1_node31_MUX_bit_math_h_l1069_c3_5488_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_iftrue := VAR_layer1_node3_MUX_bit_math_h_l761_c3_850a_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iffalse := VAR_layer1_node4_MUX_bit_math_h_l772_c3_a071_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iftrue := VAR_layer1_node5_MUX_bit_math_h_l783_c3_9883_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iffalse := VAR_layer1_node6_MUX_bit_math_h_l794_c3_cf43_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iftrue := VAR_layer1_node7_MUX_bit_math_h_l805_c3_c99c_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iffalse := VAR_layer1_node8_MUX_bit_math_h_l816_c3_fa37_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iftrue := VAR_layer1_node9_MUX_bit_math_h_l827_c3_d6c2_return_output;
     -- layer2_node9_MUX[bit_math_h_l1185_c3_30b5] LATENCY=0
     -- Inputs
     layer2_node9_MUX_bit_math_h_l1185_c3_30b5_cond <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_cond;
     layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iftrue <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iftrue;
     layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iffalse <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_iffalse;
     -- Outputs
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output := layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output;

     -- layer2_node10_MUX[bit_math_h_l1196_c3_6142] LATENCY=0
     -- Inputs
     layer2_node10_MUX_bit_math_h_l1196_c3_6142_cond <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_cond;
     layer2_node10_MUX_bit_math_h_l1196_c3_6142_iftrue <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_iftrue;
     layer2_node10_MUX_bit_math_h_l1196_c3_6142_iffalse <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_iffalse;
     -- Outputs
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output := layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output;

     -- layer2_node11_MUX[bit_math_h_l1207_c3_17d4] LATENCY=0
     -- Inputs
     layer2_node11_MUX_bit_math_h_l1207_c3_17d4_cond <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_cond;
     layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iftrue <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iftrue;
     layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iffalse <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_iffalse;
     -- Outputs
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output := layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output;

     -- layer2_node0_MUX[bit_math_h_l1086_c3_74df] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l1086_c3_74df_cond <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_cond;
     layer2_node0_MUX_bit_math_h_l1086_c3_74df_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_iftrue;
     layer2_node0_MUX_bit_math_h_l1086_c3_74df_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output := layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output;

     -- layer2_node7_MUX[bit_math_h_l1163_c3_f8a3] LATENCY=0
     -- Inputs
     layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_cond <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_cond;
     layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iftrue <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iftrue;
     layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iffalse <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_iffalse;
     -- Outputs
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output := layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output;

     -- layer2_node14_MUX[bit_math_h_l1240_c3_0287] LATENCY=0
     -- Inputs
     layer2_node14_MUX_bit_math_h_l1240_c3_0287_cond <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_cond;
     layer2_node14_MUX_bit_math_h_l1240_c3_0287_iftrue <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_iftrue;
     layer2_node14_MUX_bit_math_h_l1240_c3_0287_iffalse <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_iffalse;
     -- Outputs
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output := layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output;

     -- layer2_node4_MUX[bit_math_h_l1130_c3_d0b7] LATENCY=0
     -- Inputs
     layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_cond <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_cond;
     layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iftrue <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iftrue;
     layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iffalse <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_iffalse;
     -- Outputs
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output := layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output;

     -- layer2_node8_MUX[bit_math_h_l1174_c3_51d4] LATENCY=0
     -- Inputs
     layer2_node8_MUX_bit_math_h_l1174_c3_51d4_cond <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_cond;
     layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iftrue <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iftrue;
     layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iffalse <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_iffalse;
     -- Outputs
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output := layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output;

     -- layer2_node6_MUX[bit_math_h_l1152_c3_403d] LATENCY=0
     -- Inputs
     layer2_node6_MUX_bit_math_h_l1152_c3_403d_cond <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_cond;
     layer2_node6_MUX_bit_math_h_l1152_c3_403d_iftrue <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_iftrue;
     layer2_node6_MUX_bit_math_h_l1152_c3_403d_iffalse <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_iffalse;
     -- Outputs
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output := layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output;

     -- layer2_node5_MUX[bit_math_h_l1141_c3_a33d] LATENCY=0
     -- Inputs
     layer2_node5_MUX_bit_math_h_l1141_c3_a33d_cond <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_cond;
     layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iftrue <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iftrue;
     layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iffalse <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_iffalse;
     -- Outputs
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output := layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output;

     -- layer2_node13_MUX[bit_math_h_l1229_c3_af85] LATENCY=0
     -- Inputs
     layer2_node13_MUX_bit_math_h_l1229_c3_af85_cond <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_cond;
     layer2_node13_MUX_bit_math_h_l1229_c3_af85_iftrue <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_iftrue;
     layer2_node13_MUX_bit_math_h_l1229_c3_af85_iffalse <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_iffalse;
     -- Outputs
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output := layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output;

     -- layer2_node3_MUX[bit_math_h_l1119_c3_1d4a] LATENCY=0
     -- Inputs
     layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_cond <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_cond;
     layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iftrue <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iftrue;
     layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iffalse <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_iffalse;
     -- Outputs
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output := layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output;

     -- layer2_node12_MUX[bit_math_h_l1218_c3_74f5] LATENCY=0
     -- Inputs
     layer2_node12_MUX_bit_math_h_l1218_c3_74f5_cond <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_cond;
     layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iftrue <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iftrue;
     layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iffalse <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_iffalse;
     -- Outputs
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output := layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output;

     -- layer2_node15_MUX[bit_math_h_l1251_c3_a113] LATENCY=0
     -- Inputs
     layer2_node15_MUX_bit_math_h_l1251_c3_a113_cond <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_cond;
     layer2_node15_MUX_bit_math_h_l1251_c3_a113_iftrue <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_iftrue;
     layer2_node15_MUX_bit_math_h_l1251_c3_a113_iffalse <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_iffalse;
     -- Outputs
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output := layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output;

     -- layer2_node1_MUX[bit_math_h_l1097_c3_4739] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l1097_c3_4739_cond <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_cond;
     layer2_node1_MUX_bit_math_h_l1097_c3_4739_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_iftrue;
     layer2_node1_MUX_bit_math_h_l1097_c3_4739_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output := layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output;

     -- layer2_node2_MUX[bit_math_h_l1108_c3_c83e] LATENCY=0
     -- Inputs
     layer2_node2_MUX_bit_math_h_l1108_c3_c83e_cond <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_cond;
     layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iftrue <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iftrue;
     layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iffalse <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_iffalse;
     -- Outputs
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output := layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iffalse := VAR_layer2_node0_MUX_bit_math_h_l1086_c3_74df_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_iffalse := VAR_layer2_node10_MUX_bit_math_h_l1196_c3_6142_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_iftrue := VAR_layer2_node11_MUX_bit_math_h_l1207_c3_17d4_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_iffalse := VAR_layer2_node12_MUX_bit_math_h_l1218_c3_74f5_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_iftrue := VAR_layer2_node13_MUX_bit_math_h_l1229_c3_af85_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iffalse := VAR_layer2_node14_MUX_bit_math_h_l1240_c3_0287_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iftrue := VAR_layer2_node15_MUX_bit_math_h_l1251_c3_a113_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iftrue := VAR_layer2_node1_MUX_bit_math_h_l1097_c3_4739_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iffalse := VAR_layer2_node2_MUX_bit_math_h_l1108_c3_c83e_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iftrue := VAR_layer2_node3_MUX_bit_math_h_l1119_c3_1d4a_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_iffalse := VAR_layer2_node4_MUX_bit_math_h_l1130_c3_d0b7_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_iftrue := VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a33d_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_iffalse := VAR_layer2_node6_MUX_bit_math_h_l1152_c3_403d_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_iftrue := VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f8a3_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iffalse := VAR_layer2_node8_MUX_bit_math_h_l1174_c3_51d4_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iftrue := VAR_layer2_node9_MUX_bit_math_h_l1185_c3_30b5_return_output;
     -- layer3_node1_MUX[bit_math_h_l1279_c3_ca08] LATENCY=0
     -- Inputs
     layer3_node1_MUX_bit_math_h_l1279_c3_ca08_cond <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_cond;
     layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iftrue <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iftrue;
     layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iffalse <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_iffalse;
     -- Outputs
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output := layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output;

     -- layer3_node2_MUX[bit_math_h_l1290_c3_581b] LATENCY=0
     -- Inputs
     layer3_node2_MUX_bit_math_h_l1290_c3_581b_cond <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_cond;
     layer3_node2_MUX_bit_math_h_l1290_c3_581b_iftrue <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_iftrue;
     layer3_node2_MUX_bit_math_h_l1290_c3_581b_iffalse <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_iffalse;
     -- Outputs
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output := layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output;

     -- layer3_node6_MUX[bit_math_h_l1334_c3_d703] LATENCY=0
     -- Inputs
     layer3_node6_MUX_bit_math_h_l1334_c3_d703_cond <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_cond;
     layer3_node6_MUX_bit_math_h_l1334_c3_d703_iftrue <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_iftrue;
     layer3_node6_MUX_bit_math_h_l1334_c3_d703_iffalse <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_iffalse;
     -- Outputs
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output := layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output;

     -- layer3_node0_MUX[bit_math_h_l1268_c3_1d33] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l1268_c3_1d33_cond <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_cond;
     layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iftrue;
     layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output := layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output;

     -- layer3_node7_MUX[bit_math_h_l1345_c3_ae83] LATENCY=0
     -- Inputs
     layer3_node7_MUX_bit_math_h_l1345_c3_ae83_cond <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_cond;
     layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iftrue <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iftrue;
     layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iffalse <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_iffalse;
     -- Outputs
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output := layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output;

     -- layer3_node5_MUX[bit_math_h_l1323_c3_8487] LATENCY=0
     -- Inputs
     layer3_node5_MUX_bit_math_h_l1323_c3_8487_cond <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_cond;
     layer3_node5_MUX_bit_math_h_l1323_c3_8487_iftrue <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_iftrue;
     layer3_node5_MUX_bit_math_h_l1323_c3_8487_iffalse <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_iffalse;
     -- Outputs
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output := layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output;

     -- layer3_node3_MUX[bit_math_h_l1301_c3_778a] LATENCY=0
     -- Inputs
     layer3_node3_MUX_bit_math_h_l1301_c3_778a_cond <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_cond;
     layer3_node3_MUX_bit_math_h_l1301_c3_778a_iftrue <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_iftrue;
     layer3_node3_MUX_bit_math_h_l1301_c3_778a_iffalse <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_iffalse;
     -- Outputs
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output := layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output;

     -- layer3_node4_MUX[bit_math_h_l1312_c3_9af8] LATENCY=0
     -- Inputs
     layer3_node4_MUX_bit_math_h_l1312_c3_9af8_cond <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_cond;
     layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iftrue <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iftrue;
     layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iffalse <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_iffalse;
     -- Outputs
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output := layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output;

     -- Submodule level 5
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_iffalse := VAR_layer3_node0_MUX_bit_math_h_l1268_c3_1d33_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_iftrue := VAR_layer3_node1_MUX_bit_math_h_l1279_c3_ca08_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iffalse := VAR_layer3_node2_MUX_bit_math_h_l1290_c3_581b_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iftrue := VAR_layer3_node3_MUX_bit_math_h_l1301_c3_778a_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_iffalse := VAR_layer3_node4_MUX_bit_math_h_l1312_c3_9af8_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_iftrue := VAR_layer3_node5_MUX_bit_math_h_l1323_c3_8487_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iffalse := VAR_layer3_node6_MUX_bit_math_h_l1334_c3_d703_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iftrue := VAR_layer3_node7_MUX_bit_math_h_l1345_c3_ae83_return_output;
     -- layer4_node2_MUX[bit_math_h_l1384_c3_2032] LATENCY=0
     -- Inputs
     layer4_node2_MUX_bit_math_h_l1384_c3_2032_cond <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_cond;
     layer4_node2_MUX_bit_math_h_l1384_c3_2032_iftrue <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_iftrue;
     layer4_node2_MUX_bit_math_h_l1384_c3_2032_iffalse <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_iffalse;
     -- Outputs
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output := layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output;

     -- layer4_node0_MUX[bit_math_h_l1362_c3_0390] LATENCY=0
     -- Inputs
     layer4_node0_MUX_bit_math_h_l1362_c3_0390_cond <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_cond;
     layer4_node0_MUX_bit_math_h_l1362_c3_0390_iftrue <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_iftrue;
     layer4_node0_MUX_bit_math_h_l1362_c3_0390_iffalse <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_iffalse;
     -- Outputs
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output := layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output;

     -- layer4_node3_MUX[bit_math_h_l1395_c3_ef44] LATENCY=0
     -- Inputs
     layer4_node3_MUX_bit_math_h_l1395_c3_ef44_cond <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_cond;
     layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iftrue <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iftrue;
     layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iffalse <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_iffalse;
     -- Outputs
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output := layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output;

     -- layer4_node1_MUX[bit_math_h_l1373_c3_27d5] LATENCY=0
     -- Inputs
     layer4_node1_MUX_bit_math_h_l1373_c3_27d5_cond <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_cond;
     layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iftrue <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iftrue;
     layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iffalse <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_iffalse;
     -- Outputs
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output := layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output;

     -- Submodule level 6
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_iffalse := VAR_layer4_node0_MUX_bit_math_h_l1362_c3_0390_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_iftrue := VAR_layer4_node1_MUX_bit_math_h_l1373_c3_27d5_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iffalse := VAR_layer4_node2_MUX_bit_math_h_l1384_c3_2032_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iftrue := VAR_layer4_node3_MUX_bit_math_h_l1395_c3_ef44_return_output;
     -- layer5_node1_MUX[bit_math_h_l1423_c3_54e8] LATENCY=0
     -- Inputs
     layer5_node1_MUX_bit_math_h_l1423_c3_54e8_cond <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_cond;
     layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iftrue <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iftrue;
     layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iffalse <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_iffalse;
     -- Outputs
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output := layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output;

     -- layer5_node0_MUX[bit_math_h_l1412_c3_1733] LATENCY=0
     -- Inputs
     layer5_node0_MUX_bit_math_h_l1412_c3_1733_cond <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_cond;
     layer5_node0_MUX_bit_math_h_l1412_c3_1733_iftrue <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_iftrue;
     layer5_node0_MUX_bit_math_h_l1412_c3_1733_iffalse <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_iffalse;
     -- Outputs
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output := layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output;

     -- Submodule level 7
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iffalse := VAR_layer5_node0_MUX_bit_math_h_l1412_c3_1733_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iftrue := VAR_layer5_node1_MUX_bit_math_h_l1423_c3_54e8_return_output;
     -- layer6_node0_MUX[bit_math_h_l1440_c3_c11f] LATENCY=0
     -- Inputs
     layer6_node0_MUX_bit_math_h_l1440_c3_c11f_cond <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_cond;
     layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iftrue <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iftrue;
     layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iffalse <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_iffalse;
     -- Outputs
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output := layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output;

     -- Submodule level 8
     VAR_return_output := VAR_layer6_node0_MUX_bit_math_h_l1440_c3_c11f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
