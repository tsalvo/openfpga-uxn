-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 0
entity read_rom_byte_uxn_rom_RAM_SP_RF_1_0CLK_de264c78 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 addr0 : in unsigned(10 downto 0);
 wd : in unsigned(7 downto 0);
 we : in unsigned(0 downto 0);
 return_output : out unsigned(7 downto 0));
end read_rom_byte_uxn_rom_RAM_SP_RF_1_0CLK_de264c78;
architecture arch of read_rom_byte_uxn_rom_RAM_SP_RF_1_0CLK_de264c78 is

  signal addr : unsigned(10 downto 0) := to_unsigned(0, 11);

  signal uxn_rom : uint8_t_2048 := (
0 => to_unsigned(160, 8),
1 => to_unsigned(1, 8),
2 => to_unsigned(14, 8),
3 => to_unsigned(128, 8),
4 => to_unsigned(32, 8),
5 => to_unsigned(55, 8),
6 => to_unsigned(224, 8),
7 => to_unsigned(0, 8),
8 => to_unsigned(0, 8),
9 => to_unsigned(96, 8),
10 => to_unsigned(7, 8),
11 => to_unsigned(56, 8),
12 => to_unsigned(98, 8),
13 => to_unsigned(0, 8),
14 => to_unsigned(224, 8),
15 => to_unsigned(0, 8),
16 => to_unsigned(0, 8),
17 => to_unsigned(96, 8),
18 => to_unsigned(4, 8),
19 => to_unsigned(157, 8),
20 => to_unsigned(34, 8),
21 => to_unsigned(98, 8),
22 => to_unsigned(0, 8),
23 => to_unsigned(0, 8),
24 => to_unsigned(129, 8),
25 => to_unsigned(129, 8),
26 => to_unsigned(129, 8),
27 => to_unsigned(129, 8),
28 => to_unsigned(129, 8),
29 => to_unsigned(129, 8),
30 => to_unsigned(129, 8),
31 => to_unsigned(127, 8),
32 => to_unsigned(0, 8),
33 => to_unsigned(3, 8),
34 => to_unsigned(6, 8),
35 => to_unsigned(9, 8),
36 => to_unsigned(12, 8),
37 => to_unsigned(15, 8),
38 => to_unsigned(18, 8),
39 => to_unsigned(21, 8),
40 => to_unsigned(24, 8),
41 => to_unsigned(28, 8),
42 => to_unsigned(31, 8),
43 => to_unsigned(34, 8),
44 => to_unsigned(37, 8),
45 => to_unsigned(40, 8),
46 => to_unsigned(43, 8),
47 => to_unsigned(46, 8),
48 => to_unsigned(48, 8),
49 => to_unsigned(51, 8),
50 => to_unsigned(54, 8),
51 => to_unsigned(57, 8),
52 => to_unsigned(60, 8),
53 => to_unsigned(63, 8),
54 => to_unsigned(65, 8),
55 => to_unsigned(68, 8),
56 => to_unsigned(71, 8),
57 => to_unsigned(73, 8),
58 => to_unsigned(76, 8),
59 => to_unsigned(78, 8),
60 => to_unsigned(81, 8),
61 => to_unsigned(83, 8),
62 => to_unsigned(85, 8),
63 => to_unsigned(88, 8),
64 => to_unsigned(90, 8),
65 => to_unsigned(92, 8),
66 => to_unsigned(94, 8),
67 => to_unsigned(96, 8),
68 => to_unsigned(98, 8),
69 => to_unsigned(100, 8),
70 => to_unsigned(102, 8),
71 => to_unsigned(104, 8),
72 => to_unsigned(106, 8),
73 => to_unsigned(108, 8),
74 => to_unsigned(109, 8),
75 => to_unsigned(111, 8),
76 => to_unsigned(112, 8),
77 => to_unsigned(114, 8),
78 => to_unsigned(115, 8),
79 => to_unsigned(117, 8),
80 => to_unsigned(118, 8),
81 => to_unsigned(119, 8),
82 => to_unsigned(120, 8),
83 => to_unsigned(121, 8),
84 => to_unsigned(122, 8),
85 => to_unsigned(123, 8),
86 => to_unsigned(124, 8),
87 => to_unsigned(124, 8),
88 => to_unsigned(125, 8),
89 => to_unsigned(126, 8),
90 => to_unsigned(126, 8),
91 => to_unsigned(127, 8),
92 => to_unsigned(127, 8),
93 => to_unsigned(127, 8),
94 => to_unsigned(127, 8),
95 => to_unsigned(127, 8),
96 => to_unsigned(128, 8),
97 => to_unsigned(128, 8),
98 => to_unsigned(156, 8),
99 => to_unsigned(8, 8),
100 => to_unsigned(128, 8),
101 => to_unsigned(255, 8),
102 => to_unsigned(26, 8),
103 => to_unsigned(4, 8),
104 => to_unsigned(108, 8),
105 => to_unsigned(36, 8),
106 => to_unsigned(160, 8),
107 => to_unsigned(128, 8),
108 => to_unsigned(0, 8),
109 => to_unsigned(188, 8),
110 => to_unsigned(40, 8),
111 => to_unsigned(128, 8),
112 => to_unsigned(255, 8),
113 => to_unsigned(26, 8),
114 => to_unsigned(6, 8),
115 => to_unsigned(38, 8),
116 => to_unsigned(37, 8),
117 => to_unsigned(62, 8),
118 => to_unsigned(37, 8),
119 => to_unsigned(3, 8),
120 => to_unsigned(128, 8),
121 => to_unsigned(15, 8),
122 => to_unsigned(28, 8),
123 => to_unsigned(63, 8),
124 => to_unsigned(62, 8),
125 => to_unsigned(108, 8),
126 => to_unsigned(103, 8),
127 => to_unsigned(224, 8),
128 => to_unsigned(0, 8),
129 => to_unsigned(2, 8),
130 => to_unsigned(121, 8),
131 => to_unsigned(239, 8),
132 => to_unsigned(21, 8),
133 => to_unsigned(2, 8),
134 => to_unsigned(160, 8),
135 => to_unsigned(1, 8),
136 => to_unsigned(32, 8),
137 => to_unsigned(212, 8),
138 => to_unsigned(79, 8),
139 => to_unsigned(128, 8),
140 => to_unsigned(64, 8),
141 => to_unsigned(28, 8),
142 => to_unsigned(32, 8),
143 => to_unsigned(0, 8),
144 => to_unsigned(8, 8),
145 => to_unsigned(212, 8),
146 => to_unsigned(79, 8),
147 => to_unsigned(96, 8),
148 => to_unsigned(255, 8),
149 => to_unsigned(202, 8),
150 => to_unsigned(64, 8),
151 => to_unsigned(0, 8),
152 => to_unsigned(9, 8),
153 => to_unsigned(212, 8),
154 => to_unsigned(79, 8),
155 => to_unsigned(96, 8),
156 => to_unsigned(255, 8),
157 => to_unsigned(194, 8),
158 => to_unsigned(160, 8),
159 => to_unsigned(255, 8),
160 => to_unsigned(255, 8),
161 => to_unsigned(62, 8),
162 => to_unsigned(160, 8),
163 => to_unsigned(0, 8),
164 => to_unsigned(63, 8),
165 => to_unsigned(60, 8),
166 => to_unsigned(56, 8),
167 => to_unsigned(20, 8),
168 => to_unsigned(96, 8),
169 => to_unsigned(255, 8),
170 => to_unsigned(181, 8),
171 => to_unsigned(212, 8),
172 => to_unsigned(79, 8),
173 => to_unsigned(128, 8),
174 => to_unsigned(128, 8),
175 => to_unsigned(28, 8),
176 => to_unsigned(32, 8),
177 => to_unsigned(0, 8),
178 => to_unsigned(6, 8),
179 => to_unsigned(160, 8),
180 => to_unsigned(0, 8),
181 => to_unsigned(1, 8),
182 => to_unsigned(64, 8),
183 => to_unsigned(0, 8),
184 => to_unsigned(3, 8),
185 => to_unsigned(160, 8),
186 => to_unsigned(255, 8),
187 => to_unsigned(255, 8),
188 => to_unsigned(58, 8),
189 => to_unsigned(64, 8),
190 => to_unsigned(0, 8),
191 => to_unsigned(3, 8),
192 => to_unsigned(160, 8),
193 => to_unsigned(0, 8),
194 => to_unsigned(0, 8),
195 => to_unsigned(3, 8),
196 => to_unsigned(96, 8),
197 => to_unsigned(255, 8),
198 => to_unsigned(153, 8),
199 => to_unsigned(98, 8),
200 => to_unsigned(108, 8),
201 => to_unsigned(103, 8),
202 => to_unsigned(224, 8),
203 => to_unsigned(0, 8),
204 => to_unsigned(2, 8),
205 => to_unsigned(121, 8),
206 => to_unsigned(239, 8),
207 => to_unsigned(21, 8),
208 => to_unsigned(2, 8),
209 => to_unsigned(212, 8),
210 => to_unsigned(79, 8),
211 => to_unsigned(96, 8),
212 => to_unsigned(255, 8),
213 => to_unsigned(138, 8),
214 => to_unsigned(160, 8),
215 => to_unsigned(0, 8),
216 => to_unsigned(64, 8),
217 => to_unsigned(56, 8),
218 => to_unsigned(96, 8),
219 => to_unsigned(255, 8),
220 => to_unsigned(161, 8),
221 => to_unsigned(64, 8),
222 => to_unsigned(0, 8),
223 => to_unsigned(3, 8),
224 => to_unsigned(160, 8),
225 => to_unsigned(0, 8),
226 => to_unsigned(0, 8),
227 => to_unsigned(3, 8),
228 => to_unsigned(96, 8),
229 => to_unsigned(255, 8),
230 => to_unsigned(121, 8),
231 => to_unsigned(98, 8),
232 => to_unsigned(108, 8),
233 => to_unsigned(103, 8),
234 => to_unsigned(224, 8),
235 => to_unsigned(0, 8),
236 => to_unsigned(22, 8),
237 => to_unsigned(121, 8),
238 => to_unsigned(239, 8),
239 => to_unsigned(160, 8),
240 => to_unsigned(0, 8),
241 => to_unsigned(20, 8),
242 => to_unsigned(56, 8),
243 => to_unsigned(53, 8),
244 => to_unsigned(239, 8),
245 => to_unsigned(160, 8),
246 => to_unsigned(0, 8),
247 => to_unsigned(18, 8),
248 => to_unsigned(56, 8),
249 => to_unsigned(53, 8),
250 => to_unsigned(239, 8),
251 => to_unsigned(160, 8),
252 => to_unsigned(0, 8),
253 => to_unsigned(16, 8),
254 => to_unsigned(56, 8),
255 => to_unsigned(53, 8),
256 => to_unsigned(239, 8),
257 => to_unsigned(160, 8),
258 => to_unsigned(0, 8),
259 => to_unsigned(14, 8),
260 => to_unsigned(56, 8),
261 => to_unsigned(53, 8),
262 => to_unsigned(239, 8),
263 => to_unsigned(160, 8),
264 => to_unsigned(0, 8),
265 => to_unsigned(12, 8),
266 => to_unsigned(56, 8),
267 => to_unsigned(21, 8),
268 => to_unsigned(2, 8),
269 => to_unsigned(239, 8),
270 => to_unsigned(160, 8),
271 => to_unsigned(0, 8),
272 => to_unsigned(16, 8),
273 => to_unsigned(56, 8),
274 => to_unsigned(52, 8),
275 => to_unsigned(239, 8),
276 => to_unsigned(160, 8),
277 => to_unsigned(0, 8),
278 => to_unsigned(20, 8),
279 => to_unsigned(56, 8),
280 => to_unsigned(52, 8),
281 => to_unsigned(57, 8),
282 => to_unsigned(239, 8),
283 => to_unsigned(160, 8),
284 => to_unsigned(0, 8),
285 => to_unsigned(10, 8),
286 => to_unsigned(56, 8),
287 => to_unsigned(53, 8),
288 => to_unsigned(239, 8),
289 => to_unsigned(160, 8),
290 => to_unsigned(0, 8),
291 => to_unsigned(14, 8),
292 => to_unsigned(56, 8),
293 => to_unsigned(52, 8),
294 => to_unsigned(239, 8),
295 => to_unsigned(160, 8),
296 => to_unsigned(0, 8),
297 => to_unsigned(18, 8),
298 => to_unsigned(56, 8),
299 => to_unsigned(52, 8),
300 => to_unsigned(57, 8),
301 => to_unsigned(239, 8),
302 => to_unsigned(160, 8),
303 => to_unsigned(0, 8),
304 => to_unsigned(8, 8),
305 => to_unsigned(56, 8),
306 => to_unsigned(53, 8),
307 => to_unsigned(160, 8),
308 => to_unsigned(0, 8),
309 => to_unsigned(1, 8),
310 => to_unsigned(239, 8),
311 => to_unsigned(160, 8),
312 => to_unsigned(0, 8),
313 => to_unsigned(6, 8),
314 => to_unsigned(56, 8),
315 => to_unsigned(53, 8),
316 => to_unsigned(239, 8),
317 => to_unsigned(160, 8),
318 => to_unsigned(0, 8),
319 => to_unsigned(8, 8),
320 => to_unsigned(56, 8),
321 => to_unsigned(52, 8),
322 => to_unsigned(160, 8),
323 => to_unsigned(128, 8),
324 => to_unsigned(0, 8),
325 => to_unsigned(62, 8),
326 => to_unsigned(160, 8),
327 => to_unsigned(128, 8),
328 => to_unsigned(0, 8),
329 => to_unsigned(43, 8),
330 => to_unsigned(128, 8),
331 => to_unsigned(0, 8),
332 => to_unsigned(8, 8),
333 => to_unsigned(32, 8),
334 => to_unsigned(0, 8),
335 => to_unsigned(25, 8),
336 => to_unsigned(160, 8),
337 => to_unsigned(255, 8),
338 => to_unsigned(255, 8),
339 => to_unsigned(239, 8),
340 => to_unsigned(160, 8),
341 => to_unsigned(0, 8),
342 => to_unsigned(6, 8),
343 => to_unsigned(56, 8),
344 => to_unsigned(53, 8),
345 => to_unsigned(160, 8),
346 => to_unsigned(0, 8),
347 => to_unsigned(0, 8),
348 => to_unsigned(239, 8),
349 => to_unsigned(160, 8),
350 => to_unsigned(0, 8),
351 => to_unsigned(8, 8),
352 => to_unsigned(56, 8),
353 => to_unsigned(52, 8),
354 => to_unsigned(57, 8),
355 => to_unsigned(239, 8),
356 => to_unsigned(160, 8),
357 => to_unsigned(0, 8),
358 => to_unsigned(8, 8),
359 => to_unsigned(56, 8),
360 => to_unsigned(53, 8),
361 => to_unsigned(239, 8),
362 => to_unsigned(160, 8),
363 => to_unsigned(0, 8),
364 => to_unsigned(8, 8),
365 => to_unsigned(56, 8),
366 => to_unsigned(52, 8),
367 => to_unsigned(128, 8),
368 => to_unsigned(16, 8),
369 => to_unsigned(63, 8),
370 => to_unsigned(239, 8),
371 => to_unsigned(160, 8),
372 => to_unsigned(0, 8),
373 => to_unsigned(10, 8),
374 => to_unsigned(56, 8),
375 => to_unsigned(52, 8),
376 => to_unsigned(57, 8),
377 => to_unsigned(239, 8),
378 => to_unsigned(160, 8),
379 => to_unsigned(0, 8),
380 => to_unsigned(4, 8),
381 => to_unsigned(56, 8),
382 => to_unsigned(53, 8),
383 => to_unsigned(239, 8),
384 => to_unsigned(160, 8),
385 => to_unsigned(0, 8),
386 => to_unsigned(18, 8),
387 => to_unsigned(56, 8),
388 => to_unsigned(52, 8),
389 => to_unsigned(239, 8),
390 => to_unsigned(33, 8),
391 => to_unsigned(33, 8),
392 => to_unsigned(53, 8),
393 => to_unsigned(239, 8),
394 => to_unsigned(160, 8),
395 => to_unsigned(0, 8),
396 => to_unsigned(20, 8),
397 => to_unsigned(56, 8),
398 => to_unsigned(52, 8),
399 => to_unsigned(239, 8),
400 => to_unsigned(53, 8),
401 => to_unsigned(239, 8),
402 => to_unsigned(52, 8),
403 => to_unsigned(160, 8),
404 => to_unsigned(128, 8),
405 => to_unsigned(0, 8),
406 => to_unsigned(62, 8),
407 => to_unsigned(239, 8),
408 => to_unsigned(160, 8),
409 => to_unsigned(0, 8),
410 => to_unsigned(16, 8),
411 => to_unsigned(56, 8),
412 => to_unsigned(52, 8),
413 => to_unsigned(160, 8),
414 => to_unsigned(128, 8),
415 => to_unsigned(0, 8),
416 => to_unsigned(62, 8),
417 => to_unsigned(42, 8),
418 => to_unsigned(128, 8),
419 => to_unsigned(0, 8),
420 => to_unsigned(4, 8),
421 => to_unsigned(128, 8),
422 => to_unsigned(1, 8),
423 => to_unsigned(30, 8),
424 => to_unsigned(160, 8),
425 => to_unsigned(0, 8),
426 => to_unsigned(0, 8),
427 => to_unsigned(40, 8),
428 => to_unsigned(32, 8),
429 => to_unsigned(0, 8),
430 => to_unsigned(106, 8),
431 => to_unsigned(239, 8),
432 => to_unsigned(52, 8),
433 => to_unsigned(128, 8),
434 => to_unsigned(40, 8),
435 => to_unsigned(55, 8),
436 => to_unsigned(239, 8),
437 => to_unsigned(33, 8),
438 => to_unsigned(33, 8),
439 => to_unsigned(52, 8),
440 => to_unsigned(128, 8),
441 => to_unsigned(42, 8),
442 => to_unsigned(55, 8),
443 => to_unsigned(239, 8),
444 => to_unsigned(160, 8),
445 => to_unsigned(0, 8),
446 => to_unsigned(12, 8),
447 => to_unsigned(56, 8),
448 => to_unsigned(20, 8),
449 => to_unsigned(128, 8),
450 => to_unsigned(46, 8),
451 => to_unsigned(23, 8),
452 => to_unsigned(160, 8),
453 => to_unsigned(128, 8),
454 => to_unsigned(0, 8),
455 => to_unsigned(239, 8),
456 => to_unsigned(160, 8),
457 => to_unsigned(0, 8),
458 => to_unsigned(4, 8),
459 => to_unsigned(56, 8),
460 => to_unsigned(52, 8),
461 => to_unsigned(160, 8),
462 => to_unsigned(128, 8),
463 => to_unsigned(0, 8),
464 => to_unsigned(62, 8),
465 => to_unsigned(43, 8),
466 => to_unsigned(32, 8),
467 => to_unsigned(0, 8),
468 => to_unsigned(21, 8),
469 => to_unsigned(239, 8),
470 => to_unsigned(160, 8),
471 => to_unsigned(0, 8),
472 => to_unsigned(4, 8),
473 => to_unsigned(56, 8),
474 => to_unsigned(180, 8),
475 => to_unsigned(239, 8),
476 => to_unsigned(160, 8),
477 => to_unsigned(0, 8),
478 => to_unsigned(8, 8),
479 => to_unsigned(56, 8),
480 => to_unsigned(52, 8),
481 => to_unsigned(128, 8),
482 => to_unsigned(16, 8),
483 => to_unsigned(63, 8),
484 => to_unsigned(56, 8),
485 => to_unsigned(36, 8),
486 => to_unsigned(53, 8),
487 => to_unsigned(64, 8),
488 => to_unsigned(0, 8),
489 => to_unsigned(38, 8),
490 => to_unsigned(239, 8),
491 => to_unsigned(33, 8),
492 => to_unsigned(33, 8),
493 => to_unsigned(180, 8),
494 => to_unsigned(239, 8),
495 => to_unsigned(160, 8),
496 => to_unsigned(0, 8),
497 => to_unsigned(6, 8),
498 => to_unsigned(56, 8),
499 => to_unsigned(52, 8),
500 => to_unsigned(56, 8),
501 => to_unsigned(36, 8),
502 => to_unsigned(53, 8),
503 => to_unsigned(239, 8),
504 => to_unsigned(160, 8),
505 => to_unsigned(0, 8),
506 => to_unsigned(4, 8),
507 => to_unsigned(56, 8),
508 => to_unsigned(180, 8),
509 => to_unsigned(239, 8),
510 => to_unsigned(160, 8),
511 => to_unsigned(0, 8),
512 => to_unsigned(8, 8),
513 => to_unsigned(56, 8),
514 => to_unsigned(52, 8),
515 => to_unsigned(239, 8),
516 => to_unsigned(160, 8),
517 => to_unsigned(0, 8),
518 => to_unsigned(10, 8),
519 => to_unsigned(56, 8),
520 => to_unsigned(52, 8),
521 => to_unsigned(57, 8),
522 => to_unsigned(128, 8),
523 => to_unsigned(16, 8),
524 => to_unsigned(63, 8),
525 => to_unsigned(56, 8),
526 => to_unsigned(36, 8),
527 => to_unsigned(53, 8),
528 => to_unsigned(239, 8),
529 => to_unsigned(180, 8),
530 => to_unsigned(161, 8),
531 => to_unsigned(37, 8),
532 => to_unsigned(53, 8),
533 => to_unsigned(34, 8),
534 => to_unsigned(64, 8),
535 => to_unsigned(255, 8),
536 => to_unsigned(120, 8),
537 => to_unsigned(160, 8),
538 => to_unsigned(0, 8),
539 => to_unsigned(0, 8),
540 => to_unsigned(98, 8),
541 => to_unsigned(108, 8),
542 => to_unsigned(103, 8),
543 => to_unsigned(224, 8),
544 => to_unsigned(0, 8),
545 => to_unsigned(22, 8),
546 => to_unsigned(121, 8),
547 => to_unsigned(239, 8),
548 => to_unsigned(160, 8),
549 => to_unsigned(0, 8),
550 => to_unsigned(20, 8),
551 => to_unsigned(56, 8),
552 => to_unsigned(53, 8),
553 => to_unsigned(239, 8),
554 => to_unsigned(160, 8),
555 => to_unsigned(0, 8),
556 => to_unsigned(18, 8),
557 => to_unsigned(56, 8),
558 => to_unsigned(53, 8),
559 => to_unsigned(239, 8),
560 => to_unsigned(160, 8),
561 => to_unsigned(0, 8),
562 => to_unsigned(16, 8),
563 => to_unsigned(56, 8),
564 => to_unsigned(53, 8),
565 => to_unsigned(239, 8),
566 => to_unsigned(160, 8),
567 => to_unsigned(0, 8),
568 => to_unsigned(14, 8),
569 => to_unsigned(56, 8),
570 => to_unsigned(53, 8),
571 => to_unsigned(239, 8),
572 => to_unsigned(160, 8),
573 => to_unsigned(0, 8),
574 => to_unsigned(12, 8),
575 => to_unsigned(56, 8),
576 => to_unsigned(21, 8),
577 => to_unsigned(2, 8),
578 => to_unsigned(239, 8),
579 => to_unsigned(160, 8),
580 => to_unsigned(0, 8),
581 => to_unsigned(16, 8),
582 => to_unsigned(56, 8),
583 => to_unsigned(52, 8),
584 => to_unsigned(239, 8),
585 => to_unsigned(160, 8),
586 => to_unsigned(0, 8),
587 => to_unsigned(20, 8),
588 => to_unsigned(56, 8),
589 => to_unsigned(52, 8),
590 => to_unsigned(57, 8),
591 => to_unsigned(239, 8),
592 => to_unsigned(160, 8),
593 => to_unsigned(0, 8),
594 => to_unsigned(10, 8),
595 => to_unsigned(56, 8),
596 => to_unsigned(53, 8),
597 => to_unsigned(239, 8),
598 => to_unsigned(160, 8),
599 => to_unsigned(0, 8),
600 => to_unsigned(14, 8),
601 => to_unsigned(56, 8),
602 => to_unsigned(52, 8),
603 => to_unsigned(239, 8),
604 => to_unsigned(160, 8),
605 => to_unsigned(0, 8),
606 => to_unsigned(18, 8),
607 => to_unsigned(56, 8),
608 => to_unsigned(52, 8),
609 => to_unsigned(57, 8),
610 => to_unsigned(239, 8),
611 => to_unsigned(160, 8),
612 => to_unsigned(0, 8),
613 => to_unsigned(8, 8),
614 => to_unsigned(56, 8),
615 => to_unsigned(53, 8),
616 => to_unsigned(160, 8),
617 => to_unsigned(0, 8),
618 => to_unsigned(1, 8),
619 => to_unsigned(239, 8),
620 => to_unsigned(160, 8),
621 => to_unsigned(0, 8),
622 => to_unsigned(6, 8),
623 => to_unsigned(56, 8),
624 => to_unsigned(53, 8),
625 => to_unsigned(239, 8),
626 => to_unsigned(160, 8),
627 => to_unsigned(0, 8),
628 => to_unsigned(10, 8),
629 => to_unsigned(56, 8),
630 => to_unsigned(52, 8),
631 => to_unsigned(160, 8),
632 => to_unsigned(128, 8),
633 => to_unsigned(0, 8),
634 => to_unsigned(62, 8),
635 => to_unsigned(160, 8),
636 => to_unsigned(128, 8),
637 => to_unsigned(0, 8),
638 => to_unsigned(43, 8),
639 => to_unsigned(128, 8),
640 => to_unsigned(0, 8),
641 => to_unsigned(8, 8),
642 => to_unsigned(32, 8),
643 => to_unsigned(0, 8),
644 => to_unsigned(25, 8),
645 => to_unsigned(160, 8),
646 => to_unsigned(255, 8),
647 => to_unsigned(255, 8),
648 => to_unsigned(239, 8),
649 => to_unsigned(160, 8),
650 => to_unsigned(0, 8),
651 => to_unsigned(6, 8),
652 => to_unsigned(56, 8),
653 => to_unsigned(53, 8),
654 => to_unsigned(160, 8),
655 => to_unsigned(0, 8),
656 => to_unsigned(0, 8),
657 => to_unsigned(239, 8),
658 => to_unsigned(160, 8),
659 => to_unsigned(0, 8),
660 => to_unsigned(10, 8),
661 => to_unsigned(56, 8),
662 => to_unsigned(52, 8),
663 => to_unsigned(57, 8),
664 => to_unsigned(239, 8),
665 => to_unsigned(160, 8),
666 => to_unsigned(0, 8),
667 => to_unsigned(10, 8),
668 => to_unsigned(56, 8),
669 => to_unsigned(53, 8),
670 => to_unsigned(239, 8),
671 => to_unsigned(160, 8),
672 => to_unsigned(0, 8),
673 => to_unsigned(10, 8),
674 => to_unsigned(56, 8),
675 => to_unsigned(52, 8),
676 => to_unsigned(128, 8),
677 => to_unsigned(16, 8),
678 => to_unsigned(63, 8),
679 => to_unsigned(239, 8),
680 => to_unsigned(160, 8),
681 => to_unsigned(0, 8),
682 => to_unsigned(8, 8),
683 => to_unsigned(56, 8),
684 => to_unsigned(52, 8),
685 => to_unsigned(57, 8),
686 => to_unsigned(239, 8),
687 => to_unsigned(160, 8),
688 => to_unsigned(0, 8),
689 => to_unsigned(4, 8),
690 => to_unsigned(56, 8),
691 => to_unsigned(53, 8),
692 => to_unsigned(239, 8),
693 => to_unsigned(160, 8),
694 => to_unsigned(0, 8),
695 => to_unsigned(20, 8),
696 => to_unsigned(56, 8),
697 => to_unsigned(52, 8),
698 => to_unsigned(239, 8),
699 => to_unsigned(33, 8),
700 => to_unsigned(33, 8),
701 => to_unsigned(53, 8),
702 => to_unsigned(239, 8),
703 => to_unsigned(160, 8),
704 => to_unsigned(0, 8),
705 => to_unsigned(18, 8),
706 => to_unsigned(56, 8),
707 => to_unsigned(52, 8),
708 => to_unsigned(239, 8),
709 => to_unsigned(53, 8),
710 => to_unsigned(239, 8),
711 => to_unsigned(52, 8),
712 => to_unsigned(160, 8),
713 => to_unsigned(128, 8),
714 => to_unsigned(0, 8),
715 => to_unsigned(62, 8),
716 => to_unsigned(239, 8),
717 => to_unsigned(160, 8),
718 => to_unsigned(0, 8),
719 => to_unsigned(14, 8),
720 => to_unsigned(56, 8),
721 => to_unsigned(52, 8),
722 => to_unsigned(160, 8),
723 => to_unsigned(128, 8),
724 => to_unsigned(0, 8),
725 => to_unsigned(62, 8),
726 => to_unsigned(42, 8),
727 => to_unsigned(128, 8),
728 => to_unsigned(0, 8),
729 => to_unsigned(4, 8),
730 => to_unsigned(128, 8),
731 => to_unsigned(1, 8),
732 => to_unsigned(30, 8),
733 => to_unsigned(160, 8),
734 => to_unsigned(0, 8),
735 => to_unsigned(0, 8),
736 => to_unsigned(40, 8),
737 => to_unsigned(32, 8),
738 => to_unsigned(0, 8),
739 => to_unsigned(106, 8),
740 => to_unsigned(239, 8),
741 => to_unsigned(33, 8),
742 => to_unsigned(33, 8),
743 => to_unsigned(52, 8),
744 => to_unsigned(128, 8),
745 => to_unsigned(40, 8),
746 => to_unsigned(55, 8),
747 => to_unsigned(239, 8),
748 => to_unsigned(52, 8),
749 => to_unsigned(128, 8),
750 => to_unsigned(42, 8),
751 => to_unsigned(55, 8),
752 => to_unsigned(239, 8),
753 => to_unsigned(160, 8),
754 => to_unsigned(0, 8),
755 => to_unsigned(12, 8),
756 => to_unsigned(56, 8),
757 => to_unsigned(20, 8),
758 => to_unsigned(128, 8),
759 => to_unsigned(46, 8),
760 => to_unsigned(23, 8),
761 => to_unsigned(160, 8),
762 => to_unsigned(128, 8),
763 => to_unsigned(0, 8),
764 => to_unsigned(239, 8),
765 => to_unsigned(160, 8),
766 => to_unsigned(0, 8),
767 => to_unsigned(4, 8),
768 => to_unsigned(56, 8),
769 => to_unsigned(52, 8),
770 => to_unsigned(160, 8),
771 => to_unsigned(128, 8),
772 => to_unsigned(0, 8),
773 => to_unsigned(62, 8),
774 => to_unsigned(43, 8),
775 => to_unsigned(32, 8),
776 => to_unsigned(0, 8),
777 => to_unsigned(21, 8),
778 => to_unsigned(239, 8),
779 => to_unsigned(160, 8),
780 => to_unsigned(0, 8),
781 => to_unsigned(4, 8),
782 => to_unsigned(56, 8),
783 => to_unsigned(180, 8),
784 => to_unsigned(239, 8),
785 => to_unsigned(160, 8),
786 => to_unsigned(0, 8),
787 => to_unsigned(10, 8),
788 => to_unsigned(56, 8),
789 => to_unsigned(52, 8),
790 => to_unsigned(128, 8),
791 => to_unsigned(16, 8),
792 => to_unsigned(63, 8),
793 => to_unsigned(56, 8),
794 => to_unsigned(36, 8),
795 => to_unsigned(53, 8),
796 => to_unsigned(64, 8),
797 => to_unsigned(0, 8),
798 => to_unsigned(38, 8),
799 => to_unsigned(239, 8),
800 => to_unsigned(33, 8),
801 => to_unsigned(33, 8),
802 => to_unsigned(180, 8),
803 => to_unsigned(239, 8),
804 => to_unsigned(160, 8),
805 => to_unsigned(0, 8),
806 => to_unsigned(6, 8),
807 => to_unsigned(56, 8),
808 => to_unsigned(52, 8),
809 => to_unsigned(56, 8),
810 => to_unsigned(36, 8),
811 => to_unsigned(53, 8),
812 => to_unsigned(239, 8),
813 => to_unsigned(160, 8),
814 => to_unsigned(0, 8),
815 => to_unsigned(4, 8),
816 => to_unsigned(56, 8),
817 => to_unsigned(180, 8),
818 => to_unsigned(239, 8),
819 => to_unsigned(160, 8),
820 => to_unsigned(0, 8),
821 => to_unsigned(10, 8),
822 => to_unsigned(56, 8),
823 => to_unsigned(52, 8),
824 => to_unsigned(239, 8),
825 => to_unsigned(160, 8),
826 => to_unsigned(0, 8),
827 => to_unsigned(8, 8),
828 => to_unsigned(56, 8),
829 => to_unsigned(52, 8),
830 => to_unsigned(57, 8),
831 => to_unsigned(128, 8),
832 => to_unsigned(16, 8),
833 => to_unsigned(63, 8),
834 => to_unsigned(56, 8),
835 => to_unsigned(36, 8),
836 => to_unsigned(53, 8),
837 => to_unsigned(239, 8),
838 => to_unsigned(180, 8),
839 => to_unsigned(161, 8),
840 => to_unsigned(37, 8),
841 => to_unsigned(53, 8),
842 => to_unsigned(34, 8),
843 => to_unsigned(64, 8),
844 => to_unsigned(255, 8),
845 => to_unsigned(120, 8),
846 => to_unsigned(160, 8),
847 => to_unsigned(0, 8),
848 => to_unsigned(0, 8),
849 => to_unsigned(98, 8),
850 => to_unsigned(108, 8),
851 => to_unsigned(103, 8),
852 => to_unsigned(224, 8),
853 => to_unsigned(0, 8),
854 => to_unsigned(14, 8),
855 => to_unsigned(121, 8),
856 => to_unsigned(239, 8),
857 => to_unsigned(160, 8),
858 => to_unsigned(0, 8),
859 => to_unsigned(12, 8),
860 => to_unsigned(56, 8),
861 => to_unsigned(53, 8),
862 => to_unsigned(239, 8),
863 => to_unsigned(160, 8),
864 => to_unsigned(0, 8),
865 => to_unsigned(10, 8),
866 => to_unsigned(56, 8),
867 => to_unsigned(53, 8),
868 => to_unsigned(239, 8),
869 => to_unsigned(160, 8),
870 => to_unsigned(0, 8),
871 => to_unsigned(8, 8),
872 => to_unsigned(56, 8),
873 => to_unsigned(53, 8),
874 => to_unsigned(239, 8),
875 => to_unsigned(160, 8),
876 => to_unsigned(0, 8),
877 => to_unsigned(6, 8),
878 => to_unsigned(56, 8),
879 => to_unsigned(53, 8),
880 => to_unsigned(239, 8),
881 => to_unsigned(160, 8),
882 => to_unsigned(0, 8),
883 => to_unsigned(4, 8),
884 => to_unsigned(56, 8),
885 => to_unsigned(21, 8),
886 => to_unsigned(2, 8),
887 => to_unsigned(239, 8),
888 => to_unsigned(160, 8),
889 => to_unsigned(0, 8),
890 => to_unsigned(6, 8),
891 => to_unsigned(56, 8),
892 => to_unsigned(52, 8),
893 => to_unsigned(239, 8),
894 => to_unsigned(160, 8),
895 => to_unsigned(0, 8),
896 => to_unsigned(10, 8),
897 => to_unsigned(56, 8),
898 => to_unsigned(52, 8),
899 => to_unsigned(57, 8),
900 => to_unsigned(239, 8),
901 => to_unsigned(33, 8),
902 => to_unsigned(33, 8),
903 => to_unsigned(53, 8),
904 => to_unsigned(239, 8),
905 => to_unsigned(33, 8),
906 => to_unsigned(33, 8),
907 => to_unsigned(52, 8),
908 => to_unsigned(160, 8),
909 => to_unsigned(128, 8),
910 => to_unsigned(0, 8),
911 => to_unsigned(62, 8),
912 => to_unsigned(160, 8),
913 => to_unsigned(128, 8),
914 => to_unsigned(0, 8),
915 => to_unsigned(43, 8),
916 => to_unsigned(128, 8),
917 => to_unsigned(0, 8),
918 => to_unsigned(8, 8),
919 => to_unsigned(32, 8),
920 => to_unsigned(0, 8),
921 => to_unsigned(12, 8),
922 => to_unsigned(160, 8),
923 => to_unsigned(0, 8),
924 => to_unsigned(0, 8),
925 => to_unsigned(239, 8),
926 => to_unsigned(33, 8),
927 => to_unsigned(33, 8),
928 => to_unsigned(52, 8),
929 => to_unsigned(57, 8),
930 => to_unsigned(239, 8),
931 => to_unsigned(33, 8),
932 => to_unsigned(33, 8),
933 => to_unsigned(53, 8),
934 => to_unsigned(239, 8),
935 => to_unsigned(160, 8),
936 => to_unsigned(0, 8),
937 => to_unsigned(8, 8),
938 => to_unsigned(56, 8),
939 => to_unsigned(52, 8),
940 => to_unsigned(239, 8),
941 => to_unsigned(160, 8),
942 => to_unsigned(0, 8),
943 => to_unsigned(12, 8),
944 => to_unsigned(56, 8),
945 => to_unsigned(52, 8),
946 => to_unsigned(57, 8),
947 => to_unsigned(239, 8),
948 => to_unsigned(53, 8),
949 => to_unsigned(239, 8),
950 => to_unsigned(52, 8),
951 => to_unsigned(160, 8),
952 => to_unsigned(128, 8),
953 => to_unsigned(0, 8),
954 => to_unsigned(62, 8),
955 => to_unsigned(160, 8),
956 => to_unsigned(128, 8),
957 => to_unsigned(0, 8),
958 => to_unsigned(43, 8),
959 => to_unsigned(128, 8),
960 => to_unsigned(0, 8),
961 => to_unsigned(8, 8),
962 => to_unsigned(32, 8),
963 => to_unsigned(0, 8),
964 => to_unsigned(8, 8),
965 => to_unsigned(160, 8),
966 => to_unsigned(0, 8),
967 => to_unsigned(0, 8),
968 => to_unsigned(239, 8),
969 => to_unsigned(52, 8),
970 => to_unsigned(57, 8),
971 => to_unsigned(239, 8),
972 => to_unsigned(53, 8),
973 => to_unsigned(239, 8),
974 => to_unsigned(33, 8),
975 => to_unsigned(33, 8),
976 => to_unsigned(52, 8),
977 => to_unsigned(160, 8),
978 => to_unsigned(128, 8),
979 => to_unsigned(0, 8),
980 => to_unsigned(62, 8),
981 => to_unsigned(239, 8),
982 => to_unsigned(52, 8),
983 => to_unsigned(160, 8),
984 => to_unsigned(128, 8),
985 => to_unsigned(0, 8),
986 => to_unsigned(62, 8),
987 => to_unsigned(43, 8),
988 => to_unsigned(32, 8),
989 => to_unsigned(0, 8),
990 => to_unsigned(104, 8),
991 => to_unsigned(239, 8),
992 => to_unsigned(160, 8),
993 => to_unsigned(0, 8),
994 => to_unsigned(6, 8),
995 => to_unsigned(56, 8),
996 => to_unsigned(52, 8),
997 => to_unsigned(160, 8),
998 => to_unsigned(128, 8),
999 => to_unsigned(0, 8),
1000 => to_unsigned(62, 8),
1001 => to_unsigned(239, 8),
1002 => to_unsigned(160, 8),
1003 => to_unsigned(0, 8),
1004 => to_unsigned(10, 8),
1005 => to_unsigned(56, 8),
1006 => to_unsigned(52, 8),
1007 => to_unsigned(160, 8),
1008 => to_unsigned(128, 8),
1009 => to_unsigned(0, 8),
1010 => to_unsigned(62, 8),
1011 => to_unsigned(43, 8),
1012 => to_unsigned(32, 8),
1013 => to_unsigned(0, 8),
1014 => to_unsigned(40, 8),
1015 => to_unsigned(239, 8),
1016 => to_unsigned(160, 8),
1017 => to_unsigned(0, 8),
1018 => to_unsigned(4, 8),
1019 => to_unsigned(56, 8),
1020 => to_unsigned(20, 8),
1021 => to_unsigned(96, 8),
1022 => to_unsigned(252, 8),
1023 => to_unsigned(96, 8),
1024 => to_unsigned(239, 8),
1025 => to_unsigned(160, 8),
1026 => to_unsigned(0, 8),
1027 => to_unsigned(6, 8),
1028 => to_unsigned(56, 8),
1029 => to_unsigned(52, 8),
1030 => to_unsigned(239, 8),
1031 => to_unsigned(160, 8),
1032 => to_unsigned(0, 8),
1033 => to_unsigned(8, 8),
1034 => to_unsigned(56, 8),
1035 => to_unsigned(52, 8),
1036 => to_unsigned(239, 8),
1037 => to_unsigned(160, 8),
1038 => to_unsigned(0, 8),
1039 => to_unsigned(10, 8),
1040 => to_unsigned(56, 8),
1041 => to_unsigned(52, 8),
1042 => to_unsigned(239, 8),
1043 => to_unsigned(160, 8),
1044 => to_unsigned(0, 8),
1045 => to_unsigned(12, 8),
1046 => to_unsigned(56, 8),
1047 => to_unsigned(52, 8),
1048 => to_unsigned(96, 8),
1049 => to_unsigned(254, 8),
1050 => to_unsigned(3, 8),
1051 => to_unsigned(34, 8),
1052 => to_unsigned(64, 8),
1053 => to_unsigned(0, 8),
1054 => to_unsigned(37, 8),
1055 => to_unsigned(239, 8),
1056 => to_unsigned(160, 8),
1057 => to_unsigned(0, 8),
1058 => to_unsigned(4, 8),
1059 => to_unsigned(56, 8),
1060 => to_unsigned(20, 8),
1061 => to_unsigned(96, 8),
1062 => to_unsigned(252, 8),
1063 => to_unsigned(56, 8),
1064 => to_unsigned(239, 8),
1065 => to_unsigned(160, 8),
1066 => to_unsigned(0, 8),
1067 => to_unsigned(10, 8),
1068 => to_unsigned(56, 8),
1069 => to_unsigned(52, 8),
1070 => to_unsigned(239, 8),
1071 => to_unsigned(160, 8),
1072 => to_unsigned(0, 8),
1073 => to_unsigned(12, 8),
1074 => to_unsigned(56, 8),
1075 => to_unsigned(52, 8),
1076 => to_unsigned(239, 8),
1077 => to_unsigned(160, 8),
1078 => to_unsigned(0, 8),
1079 => to_unsigned(6, 8),
1080 => to_unsigned(56, 8),
1081 => to_unsigned(52, 8),
1082 => to_unsigned(239, 8),
1083 => to_unsigned(160, 8),
1084 => to_unsigned(0, 8),
1085 => to_unsigned(8, 8),
1086 => to_unsigned(56, 8),
1087 => to_unsigned(52, 8),
1088 => to_unsigned(96, 8),
1089 => to_unsigned(253, 8),
1090 => to_unsigned(219, 8),
1091 => to_unsigned(34, 8),
1092 => to_unsigned(64, 8),
1093 => to_unsigned(0, 8),
1094 => to_unsigned(101, 8),
1095 => to_unsigned(239, 8),
1096 => to_unsigned(160, 8),
1097 => to_unsigned(0, 8),
1098 => to_unsigned(8, 8),
1099 => to_unsigned(56, 8),
1100 => to_unsigned(52, 8),
1101 => to_unsigned(160, 8),
1102 => to_unsigned(128, 8),
1103 => to_unsigned(0, 8),
1104 => to_unsigned(62, 8),
1105 => to_unsigned(239, 8),
1106 => to_unsigned(160, 8),
1107 => to_unsigned(0, 8),
1108 => to_unsigned(12, 8),
1109 => to_unsigned(56, 8),
1110 => to_unsigned(52, 8),
1111 => to_unsigned(160, 8),
1112 => to_unsigned(128, 8),
1113 => to_unsigned(0, 8),
1114 => to_unsigned(62, 8),
1115 => to_unsigned(43, 8),
1116 => to_unsigned(32, 8),
1117 => to_unsigned(0, 8),
1118 => to_unsigned(40, 8),
1119 => to_unsigned(239, 8),
1120 => to_unsigned(160, 8),
1121 => to_unsigned(0, 8),
1122 => to_unsigned(4, 8),
1123 => to_unsigned(56, 8),
1124 => to_unsigned(20, 8),
1125 => to_unsigned(96, 8),
1126 => to_unsigned(251, 8),
1127 => to_unsigned(248, 8),
1128 => to_unsigned(239, 8),
1129 => to_unsigned(160, 8),
1130 => to_unsigned(0, 8),
1131 => to_unsigned(6, 8),
1132 => to_unsigned(56, 8),
1133 => to_unsigned(52, 8),
1134 => to_unsigned(239, 8),
1135 => to_unsigned(160, 8),
1136 => to_unsigned(0, 8),
1137 => to_unsigned(8, 8),
1138 => to_unsigned(56, 8),
1139 => to_unsigned(52, 8),
1140 => to_unsigned(239, 8),
1141 => to_unsigned(160, 8),
1142 => to_unsigned(0, 8),
1143 => to_unsigned(10, 8),
1144 => to_unsigned(56, 8),
1145 => to_unsigned(52, 8),
1146 => to_unsigned(239, 8),
1147 => to_unsigned(160, 8),
1148 => to_unsigned(0, 8),
1149 => to_unsigned(12, 8),
1150 => to_unsigned(56, 8),
1151 => to_unsigned(52, 8),
1152 => to_unsigned(96, 8),
1153 => to_unsigned(252, 8),
1154 => to_unsigned(102, 8),
1155 => to_unsigned(34, 8),
1156 => to_unsigned(64, 8),
1157 => to_unsigned(0, 8),
1158 => to_unsigned(37, 8),
1159 => to_unsigned(239, 8),
1160 => to_unsigned(160, 8),
1161 => to_unsigned(0, 8),
1162 => to_unsigned(4, 8),
1163 => to_unsigned(56, 8),
1164 => to_unsigned(20, 8),
1165 => to_unsigned(96, 8),
1166 => to_unsigned(251, 8),
1167 => to_unsigned(208, 8),
1168 => to_unsigned(239, 8),
1169 => to_unsigned(160, 8),
1170 => to_unsigned(0, 8),
1171 => to_unsigned(10, 8),
1172 => to_unsigned(56, 8),
1173 => to_unsigned(52, 8),
1174 => to_unsigned(239, 8),
1175 => to_unsigned(160, 8),
1176 => to_unsigned(0, 8),
1177 => to_unsigned(12, 8),
1178 => to_unsigned(56, 8),
1179 => to_unsigned(52, 8),
1180 => to_unsigned(239, 8),
1181 => to_unsigned(160, 8),
1182 => to_unsigned(0, 8),
1183 => to_unsigned(6, 8),
1184 => to_unsigned(56, 8),
1185 => to_unsigned(52, 8),
1186 => to_unsigned(239, 8),
1187 => to_unsigned(160, 8),
1188 => to_unsigned(0, 8),
1189 => to_unsigned(8, 8),
1190 => to_unsigned(56, 8),
1191 => to_unsigned(52, 8),
1192 => to_unsigned(96, 8),
1193 => to_unsigned(252, 8),
1194 => to_unsigned(62, 8),
1195 => to_unsigned(34, 8),
1196 => to_unsigned(160, 8),
1197 => to_unsigned(0, 8),
1198 => to_unsigned(0, 8),
1199 => to_unsigned(98, 8),
1200 => to_unsigned(108, 8),
1201 => to_unsigned(103, 8),
1202 => to_unsigned(224, 8),
1203 => to_unsigned(0, 8),
1204 => to_unsigned(18, 8),
1205 => to_unsigned(121, 8),
1206 => to_unsigned(160, 8),
1207 => to_unsigned(1, 8),
1208 => to_unsigned(23, 8),
1209 => to_unsigned(148, 8),
1210 => to_unsigned(96, 8),
1211 => to_unsigned(251, 8),
1212 => to_unsigned(163, 8),
1213 => to_unsigned(161, 8),
1214 => to_unsigned(37, 8),
1215 => to_unsigned(21, 8),
1216 => to_unsigned(2, 8),
1217 => to_unsigned(34, 8),
1218 => to_unsigned(160, 8),
1219 => to_unsigned(0, 8),
1220 => to_unsigned(0, 8),
1221 => to_unsigned(128, 8),
1222 => to_unsigned(40, 8),
1223 => to_unsigned(55, 8),
1224 => to_unsigned(160, 8),
1225 => to_unsigned(0, 8),
1226 => to_unsigned(0, 8),
1227 => to_unsigned(128, 8),
1228 => to_unsigned(42, 8),
1229 => to_unsigned(55, 8),
1230 => to_unsigned(160, 8),
1231 => to_unsigned(128, 8),
1232 => to_unsigned(46, 8),
1233 => to_unsigned(23, 8),
1234 => to_unsigned(160, 8),
1235 => to_unsigned(1, 8),
1236 => to_unsigned(0, 8),
1237 => to_unsigned(4, 8),
1238 => to_unsigned(239, 8),
1239 => to_unsigned(160, 8),
1240 => to_unsigned(0, 8),
1241 => to_unsigned(16, 8),
1242 => to_unsigned(56, 8),
1243 => to_unsigned(21, 8),
1244 => to_unsigned(2, 8),
1245 => to_unsigned(160, 8),
1246 => to_unsigned(0, 8),
1247 => to_unsigned(0, 8),
1248 => to_unsigned(239, 8),
1249 => to_unsigned(160, 8),
1250 => to_unsigned(0, 8),
1251 => to_unsigned(10, 8),
1252 => to_unsigned(56, 8),
1253 => to_unsigned(53, 8),
1254 => to_unsigned(239, 8),
1255 => to_unsigned(160, 8),
1256 => to_unsigned(0, 8),
1257 => to_unsigned(10, 8),
1258 => to_unsigned(56, 8),
1259 => to_unsigned(52, 8),
1260 => to_unsigned(160, 8),
1261 => to_unsigned(0, 8),
1262 => to_unsigned(11, 8),
1263 => to_unsigned(43, 8),
1264 => to_unsigned(128, 8),
1265 => to_unsigned(0, 8),
1266 => to_unsigned(8, 8),
1267 => to_unsigned(32, 8),
1268 => to_unsigned(1, 8),
1269 => to_unsigned(107, 8),
1270 => to_unsigned(160, 8),
1271 => to_unsigned(1, 8),
1272 => to_unsigned(23, 8),
1273 => to_unsigned(20, 8),
1274 => to_unsigned(96, 8),
1275 => to_unsigned(251, 8),
1276 => to_unsigned(99, 8),
1277 => to_unsigned(239, 8),
1278 => to_unsigned(160, 8),
1279 => to_unsigned(0, 8),
1280 => to_unsigned(10, 8),
1281 => to_unsigned(56, 8),
1282 => to_unsigned(52, 8),
1283 => to_unsigned(160, 8),
1284 => to_unsigned(0, 8),
1285 => to_unsigned(10, 8),
1286 => to_unsigned(39, 8),
1287 => to_unsigned(39, 8),
1288 => to_unsigned(59, 8),
1289 => to_unsigned(58, 8),
1290 => to_unsigned(57, 8),
1291 => to_unsigned(128, 8),
1292 => to_unsigned(128, 8),
1293 => to_unsigned(63, 8),
1294 => to_unsigned(160, 8),
1295 => to_unsigned(0, 8),
1296 => to_unsigned(10, 8),
1297 => to_unsigned(59, 8),
1298 => to_unsigned(56, 8),
1299 => to_unsigned(239, 8),
1300 => to_unsigned(160, 8),
1301 => to_unsigned(0, 8),
1302 => to_unsigned(8, 8),
1303 => to_unsigned(56, 8),
1304 => to_unsigned(21, 8),
1305 => to_unsigned(2, 8),
1306 => to_unsigned(239, 8),
1307 => to_unsigned(160, 8),
1308 => to_unsigned(0, 8),
1309 => to_unsigned(8, 8),
1310 => to_unsigned(56, 8),
1311 => to_unsigned(20, 8),
1312 => to_unsigned(128, 8),
1313 => to_unsigned(0, 8),
1314 => to_unsigned(4, 8),
1315 => to_unsigned(96, 8),
1316 => to_unsigned(251, 8),
1317 => to_unsigned(88, 8),
1318 => to_unsigned(239, 8),
1319 => to_unsigned(160, 8),
1320 => to_unsigned(0, 8),
1321 => to_unsigned(10, 8),
1322 => to_unsigned(56, 8),
1323 => to_unsigned(52, 8),
1324 => to_unsigned(160, 8),
1325 => to_unsigned(0, 8),
1326 => to_unsigned(1, 8),
1327 => to_unsigned(60, 8),
1328 => to_unsigned(96, 8),
1329 => to_unsigned(251, 8),
1330 => to_unsigned(54, 8),
1331 => to_unsigned(239, 8),
1332 => to_unsigned(160, 8),
1333 => to_unsigned(0, 8),
1334 => to_unsigned(6, 8),
1335 => to_unsigned(56, 8),
1336 => to_unsigned(53, 8),
1337 => to_unsigned(239, 8),
1338 => to_unsigned(160, 8),
1339 => to_unsigned(0, 8),
1340 => to_unsigned(8, 8),
1341 => to_unsigned(56, 8),
1342 => to_unsigned(20, 8),
1343 => to_unsigned(128, 8),
1344 => to_unsigned(0, 8),
1345 => to_unsigned(4, 8),
1346 => to_unsigned(96, 8),
1347 => to_unsigned(251, 8),
1348 => to_unsigned(132, 8),
1349 => to_unsigned(239, 8),
1350 => to_unsigned(160, 8),
1351 => to_unsigned(0, 8),
1352 => to_unsigned(10, 8),
1353 => to_unsigned(56, 8),
1354 => to_unsigned(52, 8),
1355 => to_unsigned(160, 8),
1356 => to_unsigned(0, 8),
1357 => to_unsigned(1, 8),
1358 => to_unsigned(60, 8),
1359 => to_unsigned(96, 8),
1360 => to_unsigned(251, 8),
1361 => to_unsigned(23, 8),
1362 => to_unsigned(239, 8),
1363 => to_unsigned(160, 8),
1364 => to_unsigned(0, 8),
1365 => to_unsigned(4, 8),
1366 => to_unsigned(56, 8),
1367 => to_unsigned(53, 8),
1368 => to_unsigned(239, 8),
1369 => to_unsigned(160, 8),
1370 => to_unsigned(0, 8),
1371 => to_unsigned(16, 8),
1372 => to_unsigned(56, 8),
1373 => to_unsigned(20, 8),
1374 => to_unsigned(32, 8),
1375 => to_unsigned(0, 8),
1376 => to_unsigned(208, 8),
1377 => to_unsigned(160, 8),
1378 => to_unsigned(0, 8),
1379 => to_unsigned(3, 8),
1380 => to_unsigned(239, 8),
1381 => to_unsigned(160, 8),
1382 => to_unsigned(0, 8),
1383 => to_unsigned(4, 8),
1384 => to_unsigned(56, 8),
1385 => to_unsigned(52, 8),
1386 => to_unsigned(160, 8),
1387 => to_unsigned(0, 8),
1388 => to_unsigned(179, 8),
1389 => to_unsigned(56, 8),
1390 => to_unsigned(239, 8),
1391 => to_unsigned(160, 8),
1392 => to_unsigned(0, 8),
1393 => to_unsigned(6, 8),
1394 => to_unsigned(56, 8),
1395 => to_unsigned(52, 8),
1396 => to_unsigned(160, 8),
1397 => to_unsigned(0, 8),
1398 => to_unsigned(199, 8),
1399 => to_unsigned(56, 8),
1400 => to_unsigned(239, 8),
1401 => to_unsigned(160, 8),
1402 => to_unsigned(0, 8),
1403 => to_unsigned(12, 8),
1404 => to_unsigned(56, 8),
1405 => to_unsigned(52, 8),
1406 => to_unsigned(160, 8),
1407 => to_unsigned(0, 8),
1408 => to_unsigned(179, 8),
1409 => to_unsigned(56, 8),
1410 => to_unsigned(239, 8),
1411 => to_unsigned(160, 8),
1412 => to_unsigned(0, 8),
1413 => to_unsigned(14, 8),
1414 => to_unsigned(56, 8),
1415 => to_unsigned(52, 8),
1416 => to_unsigned(160, 8),
1417 => to_unsigned(0, 8),
1418 => to_unsigned(199, 8),
1419 => to_unsigned(56, 8),
1420 => to_unsigned(96, 8),
1421 => to_unsigned(253, 8),
1422 => to_unsigned(196, 8),
1423 => to_unsigned(34, 8),
1424 => to_unsigned(160, 8),
1425 => to_unsigned(0, 8),
1426 => to_unsigned(2, 8),
1427 => to_unsigned(239, 8),
1428 => to_unsigned(160, 8),
1429 => to_unsigned(0, 8),
1430 => to_unsigned(4, 8),
1431 => to_unsigned(56, 8),
1432 => to_unsigned(52, 8),
1433 => to_unsigned(160, 8),
1434 => to_unsigned(0, 8),
1435 => to_unsigned(3, 8),
1436 => to_unsigned(58, 8),
1437 => to_unsigned(160, 8),
1438 => to_unsigned(0, 8),
1439 => to_unsigned(2, 8),
1440 => to_unsigned(96, 8),
1441 => to_unsigned(250, 8),
1442 => to_unsigned(198, 8),
1443 => to_unsigned(160, 8),
1444 => to_unsigned(0, 8),
1445 => to_unsigned(179, 8),
1446 => to_unsigned(56, 8),
1447 => to_unsigned(239, 8),
1448 => to_unsigned(160, 8),
1449 => to_unsigned(0, 8),
1450 => to_unsigned(6, 8),
1451 => to_unsigned(56, 8),
1452 => to_unsigned(52, 8),
1453 => to_unsigned(160, 8),
1454 => to_unsigned(0, 8),
1455 => to_unsigned(3, 8),
1456 => to_unsigned(58, 8),
1457 => to_unsigned(160, 8),
1458 => to_unsigned(0, 8),
1459 => to_unsigned(2, 8),
1460 => to_unsigned(96, 8),
1461 => to_unsigned(250, 8),
1462 => to_unsigned(178, 8),
1463 => to_unsigned(160, 8),
1464 => to_unsigned(0, 8),
1465 => to_unsigned(199, 8),
1466 => to_unsigned(56, 8),
1467 => to_unsigned(239, 8),
1468 => to_unsigned(160, 8),
1469 => to_unsigned(0, 8),
1470 => to_unsigned(12, 8),
1471 => to_unsigned(56, 8),
1472 => to_unsigned(52, 8),
1473 => to_unsigned(160, 8),
1474 => to_unsigned(0, 8),
1475 => to_unsigned(3, 8),
1476 => to_unsigned(58, 8),
1477 => to_unsigned(160, 8),
1478 => to_unsigned(0, 8),
1479 => to_unsigned(2, 8),
1480 => to_unsigned(96, 8),
1481 => to_unsigned(250, 8),
1482 => to_unsigned(158, 8),
1483 => to_unsigned(160, 8),
1484 => to_unsigned(0, 8),
1485 => to_unsigned(179, 8),
1486 => to_unsigned(56, 8),
1487 => to_unsigned(239, 8),
1488 => to_unsigned(160, 8),
1489 => to_unsigned(0, 8),
1490 => to_unsigned(14, 8),
1491 => to_unsigned(56, 8),
1492 => to_unsigned(52, 8),
1493 => to_unsigned(160, 8),
1494 => to_unsigned(0, 8),
1495 => to_unsigned(3, 8),
1496 => to_unsigned(58, 8),
1497 => to_unsigned(160, 8),
1498 => to_unsigned(0, 8),
1499 => to_unsigned(2, 8),
1500 => to_unsigned(96, 8),
1501 => to_unsigned(250, 8),
1502 => to_unsigned(138, 8),
1503 => to_unsigned(160, 8),
1504 => to_unsigned(0, 8),
1505 => to_unsigned(199, 8),
1506 => to_unsigned(56, 8),
1507 => to_unsigned(96, 8),
1508 => to_unsigned(253, 8),
1509 => to_unsigned(109, 8),
1510 => to_unsigned(34, 8),
1511 => to_unsigned(160, 8),
1512 => to_unsigned(0, 8),
1513 => to_unsigned(1, 8),
1514 => to_unsigned(239, 8),
1515 => to_unsigned(160, 8),
1516 => to_unsigned(0, 8),
1517 => to_unsigned(4, 8),
1518 => to_unsigned(56, 8),
1519 => to_unsigned(52, 8),
1520 => to_unsigned(160, 8),
1521 => to_unsigned(0, 8),
1522 => to_unsigned(1, 8),
1523 => to_unsigned(96, 8),
1524 => to_unsigned(250, 8),
1525 => to_unsigned(115, 8),
1526 => to_unsigned(160, 8),
1527 => to_unsigned(0, 8),
1528 => to_unsigned(179, 8),
1529 => to_unsigned(56, 8),
1530 => to_unsigned(239, 8),
1531 => to_unsigned(160, 8),
1532 => to_unsigned(0, 8),
1533 => to_unsigned(6, 8),
1534 => to_unsigned(56, 8),
1535 => to_unsigned(52, 8),
1536 => to_unsigned(160, 8),
1537 => to_unsigned(0, 8),
1538 => to_unsigned(1, 8),
1539 => to_unsigned(96, 8),
1540 => to_unsigned(250, 8),
1541 => to_unsigned(99, 8),
1542 => to_unsigned(160, 8),
1543 => to_unsigned(0, 8),
1544 => to_unsigned(199, 8),
1545 => to_unsigned(56, 8),
1546 => to_unsigned(239, 8),
1547 => to_unsigned(160, 8),
1548 => to_unsigned(0, 8),
1549 => to_unsigned(12, 8),
1550 => to_unsigned(56, 8),
1551 => to_unsigned(52, 8),
1552 => to_unsigned(160, 8),
1553 => to_unsigned(0, 8),
1554 => to_unsigned(1, 8),
1555 => to_unsigned(96, 8),
1556 => to_unsigned(250, 8),
1557 => to_unsigned(83, 8),
1558 => to_unsigned(160, 8),
1559 => to_unsigned(0, 8),
1560 => to_unsigned(179, 8),
1561 => to_unsigned(56, 8),
1562 => to_unsigned(239, 8),
1563 => to_unsigned(160, 8),
1564 => to_unsigned(0, 8),
1565 => to_unsigned(14, 8),
1566 => to_unsigned(56, 8),
1567 => to_unsigned(52, 8),
1568 => to_unsigned(160, 8),
1569 => to_unsigned(0, 8),
1570 => to_unsigned(1, 8),
1571 => to_unsigned(96, 8),
1572 => to_unsigned(250, 8),
1573 => to_unsigned(67, 8),
1574 => to_unsigned(160, 8),
1575 => to_unsigned(0, 8),
1576 => to_unsigned(199, 8),
1577 => to_unsigned(56, 8),
1578 => to_unsigned(96, 8),
1579 => to_unsigned(253, 8),
1580 => to_unsigned(38, 8),
1581 => to_unsigned(34, 8),
1582 => to_unsigned(64, 8),
1583 => to_unsigned(0, 8),
1584 => to_unsigned(11, 8),
1585 => to_unsigned(160, 8),
1586 => to_unsigned(0, 8),
1587 => to_unsigned(0, 8),
1588 => to_unsigned(4, 8),
1589 => to_unsigned(239, 8),
1590 => to_unsigned(160, 8),
1591 => to_unsigned(0, 8),
1592 => to_unsigned(16, 8),
1593 => to_unsigned(56, 8),
1594 => to_unsigned(21, 8),
1595 => to_unsigned(2, 8),
1596 => to_unsigned(239, 8),
1597 => to_unsigned(160, 8),
1598 => to_unsigned(0, 8),
1599 => to_unsigned(6, 8),
1600 => to_unsigned(56, 8),
1601 => to_unsigned(52, 8),
1602 => to_unsigned(239, 8),
1603 => to_unsigned(160, 8),
1604 => to_unsigned(0, 8),
1605 => to_unsigned(14, 8),
1606 => to_unsigned(56, 8),
1607 => to_unsigned(53, 8),
1608 => to_unsigned(239, 8),
1609 => to_unsigned(160, 8),
1610 => to_unsigned(0, 8),
1611 => to_unsigned(4, 8),
1612 => to_unsigned(56, 8),
1613 => to_unsigned(52, 8),
1614 => to_unsigned(239, 8),
1615 => to_unsigned(160, 8),
1616 => to_unsigned(0, 8),
1617 => to_unsigned(12, 8),
1618 => to_unsigned(56, 8),
1619 => to_unsigned(53, 8),
1620 => to_unsigned(239, 8),
1621 => to_unsigned(160, 8),
1622 => to_unsigned(0, 8),
1623 => to_unsigned(10, 8),
1624 => to_unsigned(56, 8),
1625 => to_unsigned(180, 8),
1626 => to_unsigned(161, 8),
1627 => to_unsigned(37, 8),
1628 => to_unsigned(53, 8),
1629 => to_unsigned(34, 8),
1630 => to_unsigned(64, 8),
1631 => to_unsigned(254, 8),
1632 => to_unsigned(133, 8),
1633 => to_unsigned(160, 8),
1634 => to_unsigned(1, 8),
1635 => to_unsigned(24, 8),
1636 => to_unsigned(128, 8),
1637 => to_unsigned(44, 8),
1638 => to_unsigned(55, 8),
1639 => to_unsigned(160, 8),
1640 => to_unsigned(0, 8),
1641 => to_unsigned(185, 8),
1642 => to_unsigned(128, 8),
1643 => to_unsigned(40, 8),
1644 => to_unsigned(55, 8),
1645 => to_unsigned(160, 8),
1646 => to_unsigned(0, 8),
1647 => to_unsigned(175, 8),
1648 => to_unsigned(128, 8),
1649 => to_unsigned(42, 8),
1650 => to_unsigned(55, 8),
1651 => to_unsigned(160, 8),
1652 => to_unsigned(1, 8),
1653 => to_unsigned(47, 8),
1654 => to_unsigned(23, 8),
1655 => to_unsigned(160, 8),
1656 => to_unsigned(1, 8),
1657 => to_unsigned(23, 8),
1658 => to_unsigned(20, 8),
1659 => to_unsigned(96, 8),
1660 => to_unsigned(249, 8),
1661 => to_unsigned(226, 8),
1662 => to_unsigned(160, 8),
1663 => to_unsigned(0, 8),
1664 => to_unsigned(32, 8),
1665 => to_unsigned(56, 8),
1666 => to_unsigned(96, 8),
1667 => to_unsigned(249, 8),
1668 => to_unsigned(249, 8),
1669 => to_unsigned(160, 8),
1670 => to_unsigned(0, 8),
1671 => to_unsigned(5, 8),
1672 => to_unsigned(96, 8),
1673 => to_unsigned(249, 8),
1674 => to_unsigned(222, 8),
1675 => to_unsigned(239, 8),
1676 => to_unsigned(33, 8),
1677 => to_unsigned(33, 8),
1678 => to_unsigned(53, 8),
1679 => to_unsigned(160, 8),
1680 => to_unsigned(1, 8),
1681 => to_unsigned(23, 8),
1682 => to_unsigned(20, 8),
1683 => to_unsigned(96, 8),
1684 => to_unsigned(249, 8),
1685 => to_unsigned(202, 8),
1686 => to_unsigned(160, 8),
1687 => to_unsigned(0, 8),
1688 => to_unsigned(32, 8),
1689 => to_unsigned(56, 8),
1690 => to_unsigned(96, 8),
1691 => to_unsigned(250, 8),
1692 => to_unsigned(44, 8),
1693 => to_unsigned(160, 8),
1694 => to_unsigned(0, 8),
1695 => to_unsigned(5, 8),
1696 => to_unsigned(96, 8),
1697 => to_unsigned(249, 8),
1698 => to_unsigned(198, 8),
1699 => to_unsigned(239, 8),
1700 => to_unsigned(53, 8),
1701 => to_unsigned(160, 8),
1702 => to_unsigned(0, 8),
1703 => to_unsigned(3, 8),
1704 => to_unsigned(239, 8),
1705 => to_unsigned(52, 8),
1706 => to_unsigned(160, 8),
1707 => to_unsigned(0, 8),
1708 => to_unsigned(179, 8),
1709 => to_unsigned(56, 8),
1710 => to_unsigned(239, 8),
1711 => to_unsigned(33, 8),
1712 => to_unsigned(33, 8),
1713 => to_unsigned(52, 8),
1714 => to_unsigned(160, 8),
1715 => to_unsigned(0, 8),
1716 => to_unsigned(199, 8),
1717 => to_unsigned(56, 8),
1718 => to_unsigned(160, 8),
1719 => to_unsigned(0, 8),
1720 => to_unsigned(179, 8),
1721 => to_unsigned(239, 8),
1722 => to_unsigned(52, 8),
1723 => to_unsigned(57, 8),
1724 => to_unsigned(160, 8),
1725 => to_unsigned(0, 8),
1726 => to_unsigned(1, 8),
1727 => to_unsigned(57, 8),
1728 => to_unsigned(160, 8),
1729 => to_unsigned(0, 8),
1730 => to_unsigned(199, 8),
1731 => to_unsigned(239, 8),
1732 => to_unsigned(33, 8),
1733 => to_unsigned(33, 8),
1734 => to_unsigned(52, 8),
1735 => to_unsigned(57, 8),
1736 => to_unsigned(160, 8),
1737 => to_unsigned(0, 8),
1738 => to_unsigned(1, 8),
1739 => to_unsigned(57, 8),
1740 => to_unsigned(96, 8),
1741 => to_unsigned(252, 8),
1742 => to_unsigned(132, 8),
1743 => to_unsigned(34, 8),
1744 => to_unsigned(160, 8),
1745 => to_unsigned(1, 8),
1746 => to_unsigned(23, 8),
1747 => to_unsigned(20, 8),
1748 => to_unsigned(96, 8),
1749 => to_unsigned(249, 8),
1750 => to_unsigned(137, 8),
1751 => to_unsigned(160, 8),
1752 => to_unsigned(0, 8),
1753 => to_unsigned(96, 8),
1754 => to_unsigned(56, 8),
1755 => to_unsigned(96, 8),
1756 => to_unsigned(249, 8),
1757 => to_unsigned(160, 8),
1758 => to_unsigned(160, 8),
1759 => to_unsigned(0, 8),
1760 => to_unsigned(5, 8),
1761 => to_unsigned(96, 8),
1762 => to_unsigned(249, 8),
1763 => to_unsigned(133, 8),
1764 => to_unsigned(239, 8),
1765 => to_unsigned(33, 8),
1766 => to_unsigned(33, 8),
1767 => to_unsigned(53, 8),
1768 => to_unsigned(160, 8),
1769 => to_unsigned(1, 8),
1770 => to_unsigned(23, 8),
1771 => to_unsigned(20, 8),
1772 => to_unsigned(96, 8),
1773 => to_unsigned(249, 8),
1774 => to_unsigned(113, 8),
1775 => to_unsigned(160, 8),
1776 => to_unsigned(0, 8),
1777 => to_unsigned(96, 8),
1778 => to_unsigned(56, 8),
1779 => to_unsigned(96, 8),
1780 => to_unsigned(249, 8),
1781 => to_unsigned(211, 8),
1782 => to_unsigned(160, 8),
1783 => to_unsigned(0, 8),
1784 => to_unsigned(5, 8),
1785 => to_unsigned(96, 8),
1786 => to_unsigned(249, 8),
1787 => to_unsigned(109, 8),
1788 => to_unsigned(239, 8),
1789 => to_unsigned(53, 8),
1790 => to_unsigned(160, 8),
1791 => to_unsigned(0, 8),
1792 => to_unsigned(3, 8),
1793 => to_unsigned(239, 8),
1794 => to_unsigned(52, 8),
1795 => to_unsigned(160, 8),
1796 => to_unsigned(0, 8),
1797 => to_unsigned(179, 8),
1798 => to_unsigned(56, 8),
1799 => to_unsigned(239, 8),
1800 => to_unsigned(33, 8),
1801 => to_unsigned(33, 8),
1802 => to_unsigned(52, 8),
1803 => to_unsigned(160, 8),
1804 => to_unsigned(0, 8),
1805 => to_unsigned(199, 8),
1806 => to_unsigned(56, 8),
1807 => to_unsigned(160, 8),
1808 => to_unsigned(0, 8),
1809 => to_unsigned(179, 8),
1810 => to_unsigned(239, 8),
1811 => to_unsigned(52, 8),
1812 => to_unsigned(57, 8),
1813 => to_unsigned(160, 8),
1814 => to_unsigned(0, 8),
1815 => to_unsigned(1, 8),
1816 => to_unsigned(57, 8),
1817 => to_unsigned(160, 8),
1818 => to_unsigned(0, 8),
1819 => to_unsigned(199, 8),
1820 => to_unsigned(239, 8),
1821 => to_unsigned(33, 8),
1822 => to_unsigned(33, 8),
1823 => to_unsigned(52, 8),
1824 => to_unsigned(57, 8),
1825 => to_unsigned(160, 8),
1826 => to_unsigned(0, 8),
1827 => to_unsigned(1, 8),
1828 => to_unsigned(57, 8),
1829 => to_unsigned(96, 8),
1830 => to_unsigned(252, 8),
1831 => to_unsigned(43, 8),
1832 => to_unsigned(34, 8),
1833 => to_unsigned(160, 8),
1834 => to_unsigned(1, 8),
1835 => to_unsigned(24, 8),
1836 => to_unsigned(128, 8),
1837 => to_unsigned(44, 8),
1838 => to_unsigned(55, 8),
1839 => to_unsigned(160, 8),
1840 => to_unsigned(0, 8),
1841 => to_unsigned(205, 8),
1842 => to_unsigned(128, 8),
1843 => to_unsigned(40, 8),
1844 => to_unsigned(55, 8),
1845 => to_unsigned(160, 8),
1846 => to_unsigned(0, 8),
1847 => to_unsigned(175, 8),
1848 => to_unsigned(128, 8),
1849 => to_unsigned(42, 8),
1850 => to_unsigned(55, 8),
1851 => to_unsigned(160, 8),
1852 => to_unsigned(49, 8),
1853 => to_unsigned(47, 8),
1854 => to_unsigned(23, 8),
1855 => to_unsigned(160, 8),
1856 => to_unsigned(0, 8),
1857 => to_unsigned(0, 8),
1858 => to_unsigned(98, 8),
1859 => to_unsigned(108, 8),
1860 => to_unsigned(103, 8),
1861 => to_unsigned(160, 8),
1862 => to_unsigned(10, 8),
1863 => to_unsigned(175, 8),
1864 => to_unsigned(128, 8),
1865 => to_unsigned(8, 8),
1866 => to_unsigned(55, 8),
1867 => to_unsigned(160, 8),
1868 => to_unsigned(15, 8),
1869 => to_unsigned(252, 8),
1870 => to_unsigned(128, 8),
1871 => to_unsigned(10, 8),
1872 => to_unsigned(55, 8),
1873 => to_unsigned(160, 8),
1874 => to_unsigned(15, 8),
1875 => to_unsigned(170, 8),
1876 => to_unsigned(128, 8),
1877 => to_unsigned(12, 8),
1878 => to_unsigned(55, 8),
1879 => to_unsigned(160, 8),
1880 => to_unsigned(1, 8),
1881 => to_unsigned(144, 8),
1882 => to_unsigned(128, 8),
1883 => to_unsigned(34, 8),
1884 => to_unsigned(55, 8),
1885 => to_unsigned(160, 8),
1886 => to_unsigned(1, 8),
1887 => to_unsigned(104, 8),
1888 => to_unsigned(128, 8),
1889 => to_unsigned(36, 8),
1890 => to_unsigned(55, 8),
1891 => to_unsigned(160, 8),
1892 => to_unsigned(0, 8),
1893 => to_unsigned(0, 8),
1894 => to_unsigned(98, 8),
1895 => to_unsigned(108, 8),
1896 => to_unsigned(0, 8),
1897 => to_unsigned(0, 8),
1898 => to_unsigned(0, 8),
1899 => to_unsigned(0, 8),
1900 => to_unsigned(0, 8),
1901 => to_unsigned(0, 8),
1902 => to_unsigned(0, 8),
1903 => to_unsigned(0, 8),
1904 => to_unsigned(0, 8),
1905 => to_unsigned(0, 8),
1906 => to_unsigned(0, 8),
1907 => to_unsigned(0, 8),
1908 => to_unsigned(0, 8),
1909 => to_unsigned(0, 8),
1910 => to_unsigned(0, 8),
1911 => to_unsigned(0, 8),
1912 => to_unsigned(0, 8),
1913 => to_unsigned(0, 8),
1914 => to_unsigned(0, 8),
1915 => to_unsigned(0, 8),
1916 => to_unsigned(0, 8),
1917 => to_unsigned(0, 8),
1918 => to_unsigned(0, 8),
1919 => to_unsigned(0, 8),
1920 => to_unsigned(0, 8),
1921 => to_unsigned(0, 8),
1922 => to_unsigned(0, 8),
1923 => to_unsigned(0, 8),
1924 => to_unsigned(0, 8),
1925 => to_unsigned(0, 8),
1926 => to_unsigned(0, 8),
1927 => to_unsigned(0, 8),
1928 => to_unsigned(0, 8),
1929 => to_unsigned(0, 8),
1930 => to_unsigned(0, 8),
1931 => to_unsigned(0, 8),
1932 => to_unsigned(0, 8),
1933 => to_unsigned(0, 8),
1934 => to_unsigned(0, 8),
1935 => to_unsigned(0, 8),
1936 => to_unsigned(0, 8),
1937 => to_unsigned(0, 8),
1938 => to_unsigned(0, 8),
1939 => to_unsigned(0, 8),
1940 => to_unsigned(0, 8),
1941 => to_unsigned(0, 8),
1942 => to_unsigned(0, 8),
1943 => to_unsigned(0, 8),
1944 => to_unsigned(0, 8),
1945 => to_unsigned(0, 8),
1946 => to_unsigned(0, 8),
1947 => to_unsigned(0, 8),
1948 => to_unsigned(0, 8),
1949 => to_unsigned(0, 8),
1950 => to_unsigned(0, 8),
1951 => to_unsigned(0, 8),
1952 => to_unsigned(0, 8),
1953 => to_unsigned(0, 8),
1954 => to_unsigned(0, 8),
1955 => to_unsigned(0, 8),
1956 => to_unsigned(0, 8),
1957 => to_unsigned(0, 8),
1958 => to_unsigned(0, 8),
1959 => to_unsigned(0, 8),
1960 => to_unsigned(0, 8),
1961 => to_unsigned(0, 8),
1962 => to_unsigned(0, 8),
1963 => to_unsigned(0, 8),
1964 => to_unsigned(0, 8),
1965 => to_unsigned(0, 8),
1966 => to_unsigned(0, 8),
1967 => to_unsigned(0, 8),
1968 => to_unsigned(0, 8),
1969 => to_unsigned(0, 8),
1970 => to_unsigned(0, 8),
1971 => to_unsigned(0, 8),
1972 => to_unsigned(0, 8),
1973 => to_unsigned(0, 8),
1974 => to_unsigned(0, 8),
1975 => to_unsigned(0, 8),
1976 => to_unsigned(0, 8),
1977 => to_unsigned(0, 8),
1978 => to_unsigned(0, 8),
1979 => to_unsigned(0, 8),
1980 => to_unsigned(0, 8),
1981 => to_unsigned(0, 8),
1982 => to_unsigned(0, 8),
1983 => to_unsigned(0, 8),
1984 => to_unsigned(0, 8),
1985 => to_unsigned(0, 8),
1986 => to_unsigned(0, 8),
1987 => to_unsigned(0, 8),
1988 => to_unsigned(0, 8),
1989 => to_unsigned(0, 8),
1990 => to_unsigned(0, 8),
1991 => to_unsigned(0, 8),
1992 => to_unsigned(0, 8),
1993 => to_unsigned(0, 8),
1994 => to_unsigned(0, 8),
1995 => to_unsigned(0, 8),
1996 => to_unsigned(0, 8),
1997 => to_unsigned(0, 8),
1998 => to_unsigned(0, 8),
1999 => to_unsigned(0, 8),
2000 => to_unsigned(0, 8),
2001 => to_unsigned(0, 8),
2002 => to_unsigned(0, 8),
2003 => to_unsigned(0, 8),
2004 => to_unsigned(0, 8),
2005 => to_unsigned(0, 8),
2006 => to_unsigned(0, 8),
2007 => to_unsigned(0, 8),
2008 => to_unsigned(0, 8),
2009 => to_unsigned(0, 8),
2010 => to_unsigned(0, 8),
2011 => to_unsigned(0, 8),
2012 => to_unsigned(0, 8),
2013 => to_unsigned(0, 8),
2014 => to_unsigned(0, 8),
2015 => to_unsigned(0, 8),
2016 => to_unsigned(0, 8),
2017 => to_unsigned(0, 8),
2018 => to_unsigned(0, 8),
2019 => to_unsigned(0, 8),
2020 => to_unsigned(0, 8),
2021 => to_unsigned(0, 8),
2022 => to_unsigned(0, 8),
2023 => to_unsigned(0, 8),
2024 => to_unsigned(0, 8),
2025 => to_unsigned(0, 8),
2026 => to_unsigned(0, 8),
2027 => to_unsigned(0, 8),
2028 => to_unsigned(0, 8),
2029 => to_unsigned(0, 8),
2030 => to_unsigned(0, 8),
2031 => to_unsigned(0, 8),
2032 => to_unsigned(0, 8),
2033 => to_unsigned(0, 8),
2034 => to_unsigned(0, 8),
2035 => to_unsigned(0, 8),
2036 => to_unsigned(0, 8),
2037 => to_unsigned(0, 8),
2038 => to_unsigned(0, 8),
2039 => to_unsigned(0, 8),
2040 => to_unsigned(0, 8),
2041 => to_unsigned(0, 8),
2042 => to_unsigned(0, 8),
2043 => to_unsigned(0, 8),
2044 => to_unsigned(0, 8),
2045 => to_unsigned(0, 8),
2046 => to_unsigned(0, 8),
2047 => to_unsigned(0, 8),
others => to_unsigned(0, 8))
;

    signal return_output_r : unsigned(7 downto 0) := to_unsigned(0, 8);
begin


addr <= addr0 ;

      process(clk) is
      begin
        if rising_edge(clk) then
          if CLOCK_ENABLE(0)='1' then            
            -- Read first
            return_output_r <= uxn_rom(to_integer(addr));
            -- RAM logic    
            if we(0) = '1' then
              uxn_rom(to_integer(addr)) <= wd; 
            end if;
          end if;
        end if;
      end process;
      -- Tie output reg to output
      return_output <= return_output_r;
      
end arch;
