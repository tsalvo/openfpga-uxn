-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity add_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end add_0CLK_f62d646e;
architecture arch of add_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l854_c6_9d7a]
signal BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l854_c1_797b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l854_c2_285d]
signal n8_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l854_c2_285d]
signal t8_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l854_c2_285d]
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l854_c2_285d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l854_c2_285d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l854_c2_285d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l854_c2_285d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l854_c2_285d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l855_c3_ddf2[uxn_opcodes_h_l855_c3_ddf2]
signal printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l859_c11_d6b2]
signal BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal n8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal t8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l859_c7_2c9a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l862_c11_93ac]
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l862_c7_2227]
signal n8_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l862_c7_2227]
signal t8_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l862_c7_2227]
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l862_c7_2227]
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l862_c7_2227]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l862_c7_2227]
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l862_c7_2227]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l862_c7_2227]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l866_c11_5987]
signal BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l866_c7_7947]
signal n8_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l866_c7_7947]
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l866_c7_7947]
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l866_c7_7947]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l866_c7_7947]
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l866_c7_7947]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l866_c7_7947]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l869_c11_ed13]
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l869_c7_e035]
signal n8_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l869_c7_e035]
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l869_c7_e035]
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c7_e035]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l869_c7_e035]
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c7_e035]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c7_e035]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l872_c30_460b]
signal sp_relative_shift_uxn_opcodes_h_l872_c30_460b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l872_c30_460b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l872_c30_460b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l875_c21_b54e]
signal BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l877_c11_d2bd]
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l877_c7_f228]
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c7_f228]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l877_c7_f228]
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a
BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_left,
BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_right,
BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output);

-- n8_MUX_uxn_opcodes_h_l854_c2_285d
n8_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l854_c2_285d_cond,
n8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
n8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- t8_MUX_uxn_opcodes_h_l854_c2_285d
t8_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l854_c2_285d_cond,
t8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
t8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d
result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_cond,
result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

-- printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2
printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2 : entity work.printf_uxn_opcodes_h_l855_c3_ddf2_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2
BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_left,
BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_right,
BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output);

-- n8_MUX_uxn_opcodes_h_l859_c7_2c9a
n8_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- t8_MUX_uxn_opcodes_h_l859_c7_2c9a
t8_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a
result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac
BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_left,
BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_right,
BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output);

-- n8_MUX_uxn_opcodes_h_l862_c7_2227
n8_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l862_c7_2227_cond,
n8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
n8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- t8_MUX_uxn_opcodes_h_l862_c7_2227
t8_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l862_c7_2227_cond,
t8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
t8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227
result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_cond,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987
BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_left,
BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_right,
BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output);

-- n8_MUX_uxn_opcodes_h_l866_c7_7947
n8_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l866_c7_7947_cond,
n8_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
n8_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947
result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_cond,
result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13
BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_left,
BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_right,
BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output);

-- n8_MUX_uxn_opcodes_h_l869_c7_e035
n8_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l869_c7_e035_cond,
n8_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
n8_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035
result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_cond,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output);

-- sp_relative_shift_uxn_opcodes_h_l872_c30_460b
sp_relative_shift_uxn_opcodes_h_l872_c30_460b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l872_c30_460b_ins,
sp_relative_shift_uxn_opcodes_h_l872_c30_460b_x,
sp_relative_shift_uxn_opcodes_h_l872_c30_460b_y,
sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_left,
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_right,
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd
BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_left,
BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_right,
BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output,
 n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output,
 n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output,
 n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output,
 n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output,
 n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output,
 sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l856_c3_4f8a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l860_c3_c570 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l864_c3_60b1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_5877 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l875_c3_2164 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l874_c3_9d67 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l869_c7_e035_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l883_l850_DUPLICATE_3857_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l856_c3_4f8a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l856_c3_4f8a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l860_c3_c570 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l860_c3_c570;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l864_c3_60b1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l864_c3_60b1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l874_c3_9d67 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l874_c3_9d67;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_5877 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_5877;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := t8;
     -- BIN_OP_PLUS[uxn_opcodes_h_l875_c21_b54e] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_left;
     BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output := BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l862_c11_93ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l872_c30_460b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l872_c30_460b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_ins;
     sp_relative_shift_uxn_opcodes_h_l872_c30_460b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_x;
     sp_relative_shift_uxn_opcodes_h_l872_c30_460b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output := sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l854_c6_9d7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l859_c11_d6b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l869_c11_ed13] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_left;
     BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output := BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l866_c11_5987] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_left;
     BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output := BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output := result.is_sp_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l869_c7_e035_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l877_c11_d2bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_9d7a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_d6b2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_93ac_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_5987_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_ed13_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_d2bd_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l875_c3_2164 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_b54e_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_6e2b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l866_l862_l859_l877_l869_DUPLICATE_5ca9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_e56d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l866_l862_l859_l854_l877_DUPLICATE_c36c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l866_l862_l859_l854_l869_DUPLICATE_19fb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_460b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iftrue := VAR_result_u8_value_uxn_opcodes_h_l875_c3_2164;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- t8_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     t8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     t8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output := t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l854_c1_797b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c7_f228] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l877_c7_f228] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output;

     -- n8_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     n8_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     n8_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output := n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output := result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l877_c7_f228] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_797b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_n8_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_f228_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_f228_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_f228_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- t8_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output := result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- n8_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     n8_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     n8_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output := n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c7_e035] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output;

     -- printf_uxn_opcodes_h_l855_c3_ddf2[uxn_opcodes_h_l855_c3_ddf2] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l855_c3_ddf2_uxn_opcodes_h_l855_c3_ddf2_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_n8_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_e035_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- n8_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     n8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     n8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output := n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- t8_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     t8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     t8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output := t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l866_c7_7947] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output := result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_7947_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l854_c2_285d_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- n8_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l862_c7_2227] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_2227_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- n8_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     n8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     n8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output := n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l859_c7_2c9a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output := result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l854_c2_285d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_2c9a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l854_c2_285d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l883_l850_DUPLICATE_3857 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l883_l850_DUPLICATE_3857_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_285d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_285d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l883_l850_DUPLICATE_3857_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l883_l850_DUPLICATE_3857_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
