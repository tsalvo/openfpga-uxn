-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity dei_0CLK_9bcaee2f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_9bcaee2f;
architecture arch of dei_0CLK_9bcaee2f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l403_c6_ad14]
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_0c95]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l403_c2_44fc]
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : device_in_result_t;

-- t8_MUX[uxn_opcodes_h_l403_c2_44fc]
signal t8_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(7 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_44fc]
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(7 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_44fc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l419_c11_11bb]
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_b4c7]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l419_c7_0c95]
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : device_in_result_t;

-- t8_MUX[uxn_opcodes_h_l419_c7_0c95]
signal t8_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(7 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_0c95]
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_0c95]
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_0c95]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_0c95]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l419_c7_0c95]
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_0c95]
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_0c95]
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l420_c30_a0a9]
signal sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l424_c9_a383]
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l424_c9_f1fa]
signal MUX_uxn_opcodes_h_l424_c9_f1fa_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_f1fa_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_f1fa_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_f1fa_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_4a37]
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_0de3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l425_c3_0d04]
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : device_in_result_t;

-- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_0d04]
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_0d04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_0d04]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l425_c3_0d04]
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_0d04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_0d04]
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(7 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_4578]
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l426_c23_4f5c]
signal device_in_uxn_opcodes_h_l426_c23_4f5c_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_4f5c_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_4f5c_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_4f5c_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_4f5c_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_7eb9]
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_986a]
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_986a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_986a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_986a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l429_c4_986a]
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(7 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_62ed( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.device_ram_address := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_device_ram_write := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;
      base.is_stack_index_flipped := ref_toks_10;
      base.is_pc_updated := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14
BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_left,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_right,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc
device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- t8_MUX_uxn_opcodes_h_l403_c2_44fc
t8_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
t8_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
t8_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc
result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb
BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_left,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_right,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95
device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- t8_MUX_uxn_opcodes_h_l419_c7_0c95
t8_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
t8_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
t8_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95
result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output);

-- sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9
sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_ins,
sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_x,
sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_y,
sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383
BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_left,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_right,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output);

-- MUX_uxn_opcodes_h_l424_c9_f1fa
MUX_uxn_opcodes_h_l424_c9_f1fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l424_c9_f1fa_cond,
MUX_uxn_opcodes_h_l424_c9_f1fa_iftrue,
MUX_uxn_opcodes_h_l424_c9_f1fa_iffalse,
MUX_uxn_opcodes_h_l424_c9_f1fa_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_expr,
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04
device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04
result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578 : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_left,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_right,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output);

-- device_in_uxn_opcodes_h_l426_c23_4f5c
device_in_uxn_opcodes_h_l426_c23_4f5c : entity work.device_in_0CLK_c6b159da port map (
clk,
device_in_uxn_opcodes_h_l426_c23_4f5c_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l426_c23_4f5c_device_address,
device_in_uxn_opcodes_h_l426_c23_4f5c_phase,
device_in_uxn_opcodes_h_l426_c23_4f5c_previous_device_ram_read,
device_in_uxn_opcodes_h_l426_c23_4f5c_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_expr,
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_cond,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a
result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_cond,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output,
 device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output,
 sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output,
 MUX_uxn_opcodes_h_l424_c9_f1fa_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output,
 device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output,
 device_in_uxn_opcodes_h_l426_c23_4f5c_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_44fc_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_3af4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_6649 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_b432 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_ff3a_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_2855_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_3941 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_217b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_2064_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_c23e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_9faa_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_2b6d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_62ed_uxn_opcodes_h_l441_l397_DUPLICATE_8a49_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := to_unsigned(0, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_right := to_unsigned(2, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_b432 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_b432;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_3af4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_3af4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iffalse := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_6649 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_6649;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iftrue := to_unsigned(1, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iffalse := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_3941 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_3941;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := t8;
     -- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_4578] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_left;
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output := BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l419_c11_11bb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_left;
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output := BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_2b6d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_2b6d_return_output := result.is_stack_write;

     -- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_7eb9] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output := UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_9faa LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_9faa_return_output := result.stack_address_sp_offset;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_44fc_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- sp_relative_shift[uxn_opcodes_h_l420_c30_a0a9] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_ins;
     sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_x <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_x;
     sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_y <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output := sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l424_c9_a383] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_left;
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output := BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_44fc_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_c23e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_c23e_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_2064 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_2064_return_output := result.device_ram_address;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l432_c23_217b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_217b_return_output := device_in_result.dei_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l403_c6_ad14] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_left;
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output := BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l425_c8_ff3a] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_ff3a_return_output := device_in_result.is_dei_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_44fc_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_ad14_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_11bb_return_output;
     VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_a383_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_4578_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_ff3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_c23e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_c23e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_c23e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_2b6d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_2b6d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_9faa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_9faa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_9faa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_217b_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_2064_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_2064_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_2064_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_53d4_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_7eb9_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_a0a9_return_output;
     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_986a] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output := has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_4a37] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output := UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_986a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l429_c4_986a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output := result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- MUX[uxn_opcodes_h_l424_c9_f1fa] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l424_c9_f1fa_cond <= VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_cond;
     MUX_uxn_opcodes_h_l424_c9_f1fa_iftrue <= VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_iftrue;
     MUX_uxn_opcodes_h_l424_c9_f1fa_iffalse <= VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_return_output := MUX_uxn_opcodes_h_l424_c9_f1fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_986a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_986a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_device_address := VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_MUX_uxn_opcodes_h_l424_c9_f1fa_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_4a37_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_986a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_986a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_986a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_986a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_986a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_b4c7] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- t8_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     t8_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     t8_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_b4c7_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_t8_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- t8_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     t8_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     t8_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_0de3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_0de3_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;
     -- device_in[uxn_opcodes_h_l426_c23_4f5c] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l426_c23_4f5c_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l426_c23_4f5c_device_address <= VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_device_address;
     device_in_uxn_opcodes_h_l426_c23_4f5c_phase <= VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_phase;
     device_in_uxn_opcodes_h_l426_c23_4f5c_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_return_output := device_in_uxn_opcodes_h_l426_c23_4f5c_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;
     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l427_c32_2855] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_2855_return_output := VAR_device_in_uxn_opcodes_h_l426_c23_4f5c_return_output.device_ram_address;

     -- device_in_result_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_2855_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_0d04] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_0d04_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_0c95] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_0c95_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_44fc] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_62ed_uxn_opcodes_h_l441_l397_DUPLICATE_8a49 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_62ed_uxn_opcodes_h_l441_l397_DUPLICATE_8a49_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_62ed(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_44fc_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_44fc_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_62ed_uxn_opcodes_h_l441_l397_DUPLICATE_8a49_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_62ed_uxn_opcodes_h_l441_l397_DUPLICATE_8a49_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
