-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 71
entity ldz2_0CLK_d662d237 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz2_0CLK_d662d237;
architecture arch of ldz2_0CLK_d662d237 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1397_c6_e275]
signal BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1397_c1_7534]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1397_c2_7cd0]
signal result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l1398_c3_95c6[uxn_opcodes_h_l1398_c3_95c6]
signal printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1402_c11_2f02]
signal BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal t8_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1402_c7_dd95]
signal result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1405_c11_c53f]
signal BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1405_c7_0003]
signal t8_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1405_c7_0003]
signal tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1405_c7_0003]
signal result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1408_c30_3f2d]
signal sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1411_c11_1025]
signal BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1411_c7_2be9]
signal result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1413_c33_30e4]
signal BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1415_c11_fb70]
signal BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1415_c7_ad67]
signal tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1415_c7_ad67]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1415_c7_ad67]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1415_c7_ad67]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1415_c7_ad67]
signal result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l1417_c3_8af3]
signal CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1419_c11_8d65]
signal BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1419_c7_9e5c]
signal tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1419_c7_9e5c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1419_c7_9e5c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1419_c7_9e5c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1419_c7_9e5c]
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1420_c3_dade]
signal BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1425_c11_e1ac]
signal BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1425_c7_378b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1425_c7_378b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1425_c7_378b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1425_c7_378b]
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l1427_c31_2575]
signal CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1429_c11_e657]
signal BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1429_c7_df0c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1429_c7_df0c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint9_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(8 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_ff87( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.u16_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275
BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_left,
BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_right,
BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output);

-- t8_MUX_uxn_opcodes_h_l1397_c2_7cd0
t8_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0
tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0
result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

-- printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6
printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6 : entity work.printf_uxn_opcodes_h_l1398_c3_95c6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02
BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_left,
BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_right,
BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output);

-- t8_MUX_uxn_opcodes_h_l1402_c7_dd95
t8_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95
tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95
result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95
result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95
result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95
result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95
result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95
result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond,
result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f
BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_left,
BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_right,
BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output);

-- t8_MUX_uxn_opcodes_h_l1405_c7_0003
t8_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
t8_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
t8_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1405_c7_0003
tmp16_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003
result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003
result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond,
result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d
sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_ins,
sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_x,
sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_y,
sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_left,
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_right,
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9
tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9
result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9
result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond,
result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4
BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_left,
BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_right,
BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70
BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_left,
BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_right,
BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67
tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_cond,
tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue,
tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse,
tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67
result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67
result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67
result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_cond,
result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output);

-- CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3
CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_x,
CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_left,
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_right,
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c
tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond,
tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue,
tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse,
tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade
BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_left,
BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_right,
BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_left,
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_right,
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output);

-- CONST_SR_8_uxn_opcodes_h_l1427_c31_2575
CONST_SR_8_uxn_opcodes_h_l1427_c31_2575 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_x,
CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657
BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_left,
BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_right,
BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c
result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c
result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output,
 t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output,
 t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output,
 t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output,
 sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output,
 tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output,
 tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output,
 CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output,
 tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output,
 CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1399_c3_fb43 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1403_c3_e3db : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1409_c22_5167_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output : unsigned(8 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1413_c22_b9fd_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1422_c3_9402 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1423_c21_2029_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1426_c3_039b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1427_c21_52a9_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1405_l1397_l1402_DUPLICATE_518c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_7b26_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_9990_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a_return_output : unsigned(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1420_l1416_DUPLICATE_2bfd_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1434_l1392_DUPLICATE_4187_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1399_c3_fb43 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1399_c3_fb43;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1426_c3_039b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1426_c3_039b;
     VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1403_c3_e3db := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1403_c3_e3db;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1422_c3_9402 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1422_c3_9402;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := t8;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_left := tmp16;
     VAR_CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l1419_c11_8d65] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_left;
     BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output := BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1405_l1397_l1402_DUPLICATE_518c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1405_l1397_l1402_DUPLICATE_518c_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1415_c11_fb70] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_left;
     BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output := BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l1427_c31_2575] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_x <= VAR_CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output := CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1405_c11_c53f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1413_c33_30e4] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1402_c11_2f02] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_left;
     BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output := BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1429_c11_e657] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_left;
     BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output := BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1408_c30_3f2d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_ins;
     sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_x;
     sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output := sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output := result.u8_value;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1420_l1416_DUPLICATE_2bfd LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1420_l1416_DUPLICATE_2bfd_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_7b26 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_7b26_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1425_c11_e1ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1409_c22_5167] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1409_c22_5167_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1411_c11_1025] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_left;
     BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output := BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_9990 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_9990_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1397_c6_e275] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_left;
     BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output := BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1397_c6_e275_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c11_2f02_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c11_c53f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_1025_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1415_c11_fb70_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_8d65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_e1ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1429_c11_e657_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1409_c22_5167_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1420_l1416_DUPLICATE_2bfd_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1420_l1416_DUPLICATE_2bfd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1405_l1397_l1402_DUPLICATE_518c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1405_l1397_l1402_DUPLICATE_518c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1405_l1397_l1402_DUPLICATE_518c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_9990_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_9990_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_9990_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1425_l1419_l1415_l1411_DUPLICATE_251e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_7b26_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_7b26_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1397_l1411_l1402_DUPLICATE_7b26_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1405_l1402_l1429_l1397_l1425_l1415_l1411_DUPLICATE_ee99_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1415_l1405_l1411_l1425_DUPLICATE_df6a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1405_l1402_l1397_l1425_l1415_l1411_DUPLICATE_62e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1408_c30_3f2d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1429_c7_df0c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1413_c22_b9fd] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1413_c22_b9fd_return_output := CAST_TO_uint16_t_uint9_t(
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1413_c33_30e4_return_output);

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1425_c7_378b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1427_c21_52a9] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1427_c21_52a9_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l1427_c31_2575_return_output);

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1420_c3_dade] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_left;
     BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output := BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1397_c1_7534] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1429_c7_df0c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l1417_c3_8af3] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_x <= VAR_CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output := CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     t8_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     t8_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- Submodule level 2
     VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1413_c22_b9fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1427_c21_52a9_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l1417_c3_8af3_return_output;
     VAR_printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1397_c1_7534_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1429_c7_df0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1425_c7_378b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- printf_uxn_opcodes_h_l1398_c3_95c6[uxn_opcodes_h_l1398_c3_95c6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1398_c3_95c6_uxn_opcodes_h_l1398_c3_95c6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- tmp16_MUX[uxn_opcodes_h_l1419_c7_9e5c] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond;
     tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output := tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1425_c7_378b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1419_c7_9e5c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1423_c21_2029] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1423_c21_2029_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l1420_c3_dade_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1425_c7_378b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1423_c21_2029_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_378b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1419_c7_9e5c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1415_c7_ad67] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_cond;
     tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output := tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1415_c7_ad67] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1419_c7_9e5c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1419_c7_9e5c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_9e5c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1415_c7_ad67] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1415_c7_ad67] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1415_c7_ad67] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output := result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1415_c7_ad67_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1411_c7_2be9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1411_c7_2be9_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1405_c7_0003] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output := result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1405_c7_0003_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1402_c7_dd95] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;

     -- Submodule level 8
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1402_c7_dd95_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1397_c2_7cd0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1434_l1392_DUPLICATE_4187 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1434_l1392_DUPLICATE_4187_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ff87(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1397_c2_7cd0_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1434_l1392_DUPLICATE_4187_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1434_l1392_DUPLICATE_4187_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
