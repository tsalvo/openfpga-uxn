-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity equ_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_85d5529e;
architecture arch of equ_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1114_c6_1d58]
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1114_c1_39bd]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal t8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal n8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1114_c2_36ab]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l1115_c3_8226[uxn_opcodes_h_l1115_c3_8226]
signal printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1119_c11_e00e]
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1119_c7_2173]
signal t8_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1119_c7_2173]
signal n8_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1119_c7_2173]
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1119_c7_2173]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1119_c7_2173]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1119_c7_2173]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1119_c7_2173]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1119_c7_2173]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1122_c11_7f09]
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1122_c7_1ab5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1125_c11_261e]
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1125_c7_0438]
signal n8_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1125_c7_0438]
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1125_c7_0438]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1125_c7_0438]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1125_c7_0438]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1125_c7_0438]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1125_c7_0438]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1128_c30_b8c8]
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1131_c21_f22e]
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1131_c21_f4d8]
signal MUX_uxn_opcodes_h_l1131_c21_f4d8_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_f4d8_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_f4d8_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1133_c11_8e44]
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c7_a4af]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c7_a4af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c7_a4af]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_left,
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_right,
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output);

-- t8_MUX_uxn_opcodes_h_l1114_c2_36ab
t8_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- n8_MUX_uxn_opcodes_h_l1114_c2_36ab
n8_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

-- printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226
printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226 : entity work.printf_uxn_opcodes_h_l1115_c3_8226_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_left,
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_right,
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output);

-- t8_MUX_uxn_opcodes_h_l1119_c7_2173
t8_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
t8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
t8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- n8_MUX_uxn_opcodes_h_l1119_c7_2173
n8_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
n8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
n8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_left,
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_right,
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output);

-- t8_MUX_uxn_opcodes_h_l1122_c7_1ab5
t8_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- n8_MUX_uxn_opcodes_h_l1122_c7_1ab5
n8_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_left,
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_right,
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output);

-- n8_MUX_uxn_opcodes_h_l1125_c7_0438
n8_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
n8_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
n8_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8
sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_ins,
sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_x,
sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_y,
sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_left,
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_right,
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output);

-- MUX_uxn_opcodes_h_l1131_c21_f4d8
MUX_uxn_opcodes_h_l1131_c21_f4d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1131_c21_f4d8_cond,
MUX_uxn_opcodes_h_l1131_c21_f4d8_iftrue,
MUX_uxn_opcodes_h_l1131_c21_f4d8_iffalse,
MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_left,
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_right,
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output,
 t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output,
 t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output,
 t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output,
 n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output,
 sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output,
 MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_1575 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_9b3d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_bad9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_55d8_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1139_l1110_DUPLICATE_2e97_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_bad9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_bad9;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_9b3d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_9b3d;
     VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_1575 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_1575;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_55d8 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_55d8_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1128_c30_b8c8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_ins;
     sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_x;
     sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output := sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1131_c21_f22e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1125_c11_261e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1119_c11_e00e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1133_c11_8e44] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_left;
     BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output := BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1122_c11_7f09] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_left;
     BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output := BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1114_c6_1d58] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_left;
     BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output := BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_1d58_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_e00e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_7f09_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_261e_return_output;
     VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_f22e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_8e44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_96f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_47a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_70a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1119_l1133_l1122_l1114_DUPLICATE_c0ba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_55d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_55d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1125_l1119_l1122_l1114_DUPLICATE_43d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_b8c8_return_output;
     -- n8_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     n8_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     n8_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1114_c1_39bd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c7_a4af] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- MUX[uxn_opcodes_h_l1131_c21_f4d8] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1131_c21_f4d8_cond <= VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_cond;
     MUX_uxn_opcodes_h_l1131_c21_f4d8_iftrue <= VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_iftrue;
     MUX_uxn_opcodes_h_l1131_c21_f4d8_iffalse <= VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output := MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c7_a4af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c7_a4af] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output;

     -- t8_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue := VAR_MUX_uxn_opcodes_h_l1131_c21_f4d8_return_output;
     VAR_printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_39bd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_a4af_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- t8_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     t8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     t8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- n8_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- printf_uxn_opcodes_h_l1115_c3_8226[uxn_opcodes_h_l1115_c3_8226] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1115_c3_8226_uxn_opcodes_h_l1115_c3_8226_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1125_c7_0438] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0438_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- n8_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     n8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     n8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1122_c7_1ab5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- t8_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_1ab5_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- n8_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1119_c7_2173] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output := result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_2173_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1114_c2_36ab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1139_l1110_DUPLICATE_2e97 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1139_l1110_DUPLICATE_2e97_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_36ab_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1139_l1110_DUPLICATE_2e97_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1139_l1110_DUPLICATE_2e97_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
