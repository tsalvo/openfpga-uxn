-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity eor_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_f62d646e;
architecture arch of eor_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1133_c6_6e2a]
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1133_c1_3853]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1133_c2_688d]
signal n8_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1133_c2_688d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1133_c2_688d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c2_688d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c2_688d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c2_688d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1133_c2_688d]
signal result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1133_c2_688d]
signal t8_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1134_c3_2287[uxn_opcodes_h_l1134_c3_2287]
signal printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1138_c11_0276]
signal BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal n8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1138_c7_45b0]
signal t8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1141_c11_c0d1]
signal BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1141_c7_675b]
signal n8_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1141_c7_675b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1141_c7_675b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1141_c7_675b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1141_c7_675b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1141_c7_675b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1141_c7_675b]
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1141_c7_675b]
signal t8_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1145_c11_6d1c]
signal BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1145_c7_0bcd]
signal result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1148_c11_556c]
signal BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal n8_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1148_c7_f54b]
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1151_c30_258d]
signal sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1154_c21_4fff]
signal BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1156_c11_0df2]
signal BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1156_c7_d5e5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1156_c7_d5e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1156_c7_d5e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a
BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_left,
BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_right,
BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output);

-- n8_MUX_uxn_opcodes_h_l1133_c2_688d
n8_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
n8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
n8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d
result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- t8_MUX_uxn_opcodes_h_l1133_c2_688d
t8_MUX_uxn_opcodes_h_l1133_c2_688d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1133_c2_688d_cond,
t8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue,
t8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse,
t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

-- printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287
printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287 : entity work.printf_uxn_opcodes_h_l1134_c3_2287_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276
BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_left,
BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_right,
BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output);

-- n8_MUX_uxn_opcodes_h_l1138_c7_45b0
n8_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0
result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- t8_MUX_uxn_opcodes_h_l1138_c7_45b0
t8_MUX_uxn_opcodes_h_l1138_c7_45b0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond,
t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue,
t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse,
t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_left,
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_right,
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output);

-- n8_MUX_uxn_opcodes_h_l1141_c7_675b
n8_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
n8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
n8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- t8_MUX_uxn_opcodes_h_l1141_c7_675b
t8_MUX_uxn_opcodes_h_l1141_c7_675b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1141_c7_675b_cond,
t8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue,
t8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse,
t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c
BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_left,
BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_right,
BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output);

-- n8_MUX_uxn_opcodes_h_l1145_c7_0bcd
n8_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd
result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd
result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd
result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd
result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_left,
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_right,
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output);

-- n8_MUX_uxn_opcodes_h_l1148_c7_f54b
n8_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1151_c30_258d
sp_relative_shift_uxn_opcodes_h_l1151_c30_258d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_ins,
sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_x,
sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_y,
sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff
BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_left,
BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_right,
BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2
BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_left,
BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_right,
BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5
result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5
result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5
result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output,
 n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output,
 n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output,
 n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output,
 n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output,
 n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1135_c3_6738 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1139_c3_7cc1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1143_c3_803a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1146_c3_7e3a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1153_c3_2271 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1148_c7_f54b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1162_l1129_DUPLICATE_e014_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1139_c3_7cc1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1139_c3_7cc1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1146_c3_7e3a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1146_c3_7e3a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1143_c3_803a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1143_c3_803a;
     VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1153_c3_2271 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1153_c3_2271;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1135_c3_6738 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1135_c3_6738;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1138_c11_0276] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_left;
     BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output := BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1133_c6_6e2a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1156_c11_0df2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output := result.sp_relative_shift;

     -- BIN_OP_XOR[uxn_opcodes_h_l1154_c21_4fff] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_left;
     BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output := BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1148_c11_556c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1151_c30_258d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_ins;
     sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_x;
     sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output := sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1145_c11_6d1c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1148_c7_f54b_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1141_c11_c0d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c6_6e2a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c11_0276_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_c0d1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1145_c11_6d1c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_556c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1156_c11_0df2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1154_c21_4fff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_2f0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1141_l1138_l1156_l1148_l1145_DUPLICATE_8344_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_da33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1156_l1145_DUPLICATE_5997_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1141_l1138_l1133_l1148_l1145_DUPLICATE_e939_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1151_c30_258d_return_output;
     -- t8_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     t8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     t8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1156_c7_d5e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1156_c7_d5e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1133_c1_3853] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output;

     -- n8_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1156_c7_d5e5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1133_c1_3853_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1156_c7_d5e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1148_c7_f54b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;

     -- printf_uxn_opcodes_h_l1134_c3_2287[uxn_opcodes_h_l1134_c3_2287] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1134_c3_2287_uxn_opcodes_h_l1134_c3_2287_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- n8_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_f54b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     t8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     t8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1145_c7_0bcd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;

     -- n8_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     n8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     n8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1145_c7_0bcd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1141_c7_675b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_675b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- n8_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     n8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     n8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1138_c7_45b0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c7_45b0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c2_688d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1162_l1129_DUPLICATE_e014 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1162_l1129_DUPLICATE_e014_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c2_688d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1133_c2_688d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1162_l1129_DUPLICATE_e014_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1162_l1129_DUPLICATE_e014_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
