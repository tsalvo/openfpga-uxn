-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc_0CLK_3045e391 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_3045e391;
architecture arch of inc_0CLK_3045e391 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1433_c6_eb7b]
signal BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1433_c1_a084]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1433_c2_5b9b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1434_c3_1e14[uxn_opcodes_h_l1434_c3_1e14]
signal printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1438_c11_42af]
signal BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal t8_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1438_c7_cc70]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1441_c11_7391]
signal BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal t8_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1441_c7_d36f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1444_c32_580d]
signal BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1444_c32_dae5]
signal BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1444_c32_1f31]
signal MUX_uxn_opcodes_h_l1444_c32_1f31_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1444_c32_1f31_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1444_c32_1f31_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1444_c32_1f31_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1446_c11_6c55]
signal BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1446_c7_5f1c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1446_c7_5f1c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1446_c7_5f1c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1446_c7_5f1c]
signal result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1446_c7_5f1c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1450_c24_bc52]
signal BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1452_c11_3067]
signal BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1452_c7_1925]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1452_c7_1925]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_53ff( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_value := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b
BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_left,
BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_right,
BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output);

-- t8_MUX_uxn_opcodes_h_l1433_c2_5b9b
t8_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b
result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b
result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b
result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b
result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

-- printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14
printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14 : entity work.printf_uxn_opcodes_h_l1434_c3_1e14_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af
BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_left,
BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_right,
BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output);

-- t8_MUX_uxn_opcodes_h_l1438_c7_cc70
t8_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70
result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70
result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70
result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70
result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70
result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_left,
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_right,
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output);

-- t8_MUX_uxn_opcodes_h_l1441_c7_d36f
t8_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f
result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f
result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d
BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_left,
BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_right,
BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5
BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_left,
BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_right,
BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output);

-- MUX_uxn_opcodes_h_l1444_c32_1f31
MUX_uxn_opcodes_h_l1444_c32_1f31 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1444_c32_1f31_cond,
MUX_uxn_opcodes_h_l1444_c32_1f31_iftrue,
MUX_uxn_opcodes_h_l1444_c32_1f31_iffalse,
MUX_uxn_opcodes_h_l1444_c32_1f31_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55
BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_left,
BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_right,
BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c
result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c
result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c
result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond,
result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c
result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52
BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_left,
BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_right,
BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067
BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_left,
BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_right,
BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925
result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925
result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output,
 t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output,
 t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output,
 t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output,
 MUX_uxn_opcodes_h_l1444_c32_1f31_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1435_c3_b87d : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_0b54 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1449_c3_6fe7 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1450_c3_b1ad : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1441_l1433_l1438_DUPLICATE_c9ee_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1433_l1446_l1438_DUPLICATE_56bc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1441_l1446_DUPLICATE_be4b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l1457_l1429_DUPLICATE_2486_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_right := to_unsigned(128, 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_0b54 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_0b54;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_right := to_unsigned(3, 2);
     VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1449_c3_6fe7 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1449_c3_6fe7;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1435_c3_b87d := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1435_c3_b87d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1446_c11_6c55] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_left;
     BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output := BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e_return_output := result.is_opc_done;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1441_l1433_l1438_DUPLICATE_c9ee LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1441_l1433_l1438_DUPLICATE_c9ee_return_output := result.sp_relative_shift;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1450_c24_bc52] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1441_c11_7391] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_left;
     BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output := BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1433_c6_eb7b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1452_c11_3067] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_left;
     BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output := BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1441_l1446_DUPLICATE_be4b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1441_l1446_DUPLICATE_be4b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_AND[uxn_opcodes_h_l1444_c32_580d] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_left;
     BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output := BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1433_l1446_l1438_DUPLICATE_56bc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1433_l1446_l1438_DUPLICATE_56bc_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1438_c11_42af] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_left;
     BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output := BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a_return_output := result.stack_value;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1444_c32_580d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1433_c6_eb7b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1438_c11_42af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_7391_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1446_c11_6c55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1452_c11_3067_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1450_c3_b1ad := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1450_c24_bc52_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1441_l1433_l1438_DUPLICATE_c9ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1441_l1433_l1438_DUPLICATE_c9ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1441_l1433_l1438_DUPLICATE_c9ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1441_l1446_l1438_l1452_DUPLICATE_934e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1433_l1446_l1438_DUPLICATE_56bc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1433_l1446_l1438_DUPLICATE_56bc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1433_l1446_l1438_DUPLICATE_56bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1441_l1433_l1438_l1452_DUPLICATE_d802_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1441_l1446_DUPLICATE_be4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1441_l1446_DUPLICATE_be4b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1441_l1433_l1446_l1438_DUPLICATE_1e7a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1450_c3_b1ad;
     -- t8_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1433_c1_a084] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1452_c7_1925] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1446_c7_5f1c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1444_c32_dae5] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_left;
     BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output := BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1446_c7_5f1c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1446_c7_5f1c] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output := result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1452_c7_1925] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1444_c32_dae5_return_output;
     VAR_printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1433_c1_a084_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1452_c7_1925_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1452_c7_1925_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     -- printf_uxn_opcodes_h_l1434_c3_1e14[uxn_opcodes_h_l1434_c3_1e14] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1434_c3_1e14_uxn_opcodes_h_l1434_c3_1e14_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_value_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- MUX[uxn_opcodes_h_l1444_c32_1f31] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1444_c32_1f31_cond <= VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_cond;
     MUX_uxn_opcodes_h_l1444_c32_1f31_iftrue <= VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_iftrue;
     MUX_uxn_opcodes_h_l1444_c32_1f31_iffalse <= VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_return_output := MUX_uxn_opcodes_h_l1444_c32_1f31_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1446_c7_5f1c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1446_c7_5f1c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue := VAR_MUX_uxn_opcodes_h_l1444_c32_1f31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1446_c7_5f1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1441_c7_d36f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1441_c7_d36f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1438_c7_cc70] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1438_c7_cc70_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1433_c2_5b9b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l1457_l1429_DUPLICATE_2486 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l1457_l1429_DUPLICATE_2486_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_53ff(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1433_c2_5b9b_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l1457_l1429_DUPLICATE_2486_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l1457_l1429_DUPLICATE_2486_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
