-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2175_c6_b90a]
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2175_c2_7ebc]
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_a886]
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2188_c7_73c0]
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2191_c11_5df8]
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2191_c7_19b3]
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2193_c30_9d2f]
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_890c]
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2198_c7_786e]
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_786e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_786e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_786e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_786e]
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_left,
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_right,
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc
t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc
t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_left,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_right,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0
t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0
t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_left,
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_right,
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3
t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3
t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f
sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_ins,
sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_x,
sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_y,
sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_left,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_right,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2198_c7_786e
t16_low_MUX_uxn_opcodes_h_l2198_c7_786e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_cond,
t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue,
t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse,
t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output,
 t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output,
 t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output,
 t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output,
 sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output,
 t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_6dbc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_418c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_fac8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_ac83 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_97b8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_dc43 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_786e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_79a1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_0e7e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2191_l2198_l2188_DUPLICATE_a29f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2191_l2188_DUPLICATE_3ac5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2171_l2206_DUPLICATE_25ef_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_97b8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_97b8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_6dbc := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_6dbc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_418c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_418c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_fac8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_fac8;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_ac83 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_ac83;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_dc43 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_dc43;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse := t16_low;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2191_l2198_l2188_DUPLICATE_a29f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2191_l2198_l2188_DUPLICATE_a29f_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2191_c11_5df8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_890c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_79a1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_79a1_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output := result.is_stack_index_flipped;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2191_l2188_DUPLICATE_3ac5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2191_l2188_DUPLICATE_3ac5_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2193_c30_9d2f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_ins;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_x;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output := sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2175_c6_b90a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_a886] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_left;
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output := BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_0e7e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_0e7e_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2198_c7_786e] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_786e_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output := result.is_ram_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b90a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_a886_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_5df8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_890c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_0e7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_0e7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2191_l2198_l2188_DUPLICATE_a29f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2191_l2198_l2188_DUPLICATE_a29f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2191_l2198_l2188_DUPLICATE_a29f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2191_l2188_DUPLICATE_3ac5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2191_l2188_DUPLICATE_3ac5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_79a1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_79a1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_79a1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_7ebc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_786e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_9d2f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_786e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_786e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2198_c7_786e] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_cond;
     t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output := t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_786e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_786e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_786e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2191_c7_19b3] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_cond;
     t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output := t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_19b3_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_73c0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_73c0_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2175_c2_7ebc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2171_l2206_DUPLICATE_25ef LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2171_l2206_DUPLICATE_25ef_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_7ebc_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2171_l2206_DUPLICATE_25ef_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2171_l2206_DUPLICATE_25ef_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
