-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity dup2_0CLK_e4095020 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup2_0CLK_e4095020;
architecture arch of dup2_0CLK_e4095020 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2815_c6_813e]
signal BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2815_c2_1cec]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2828_c11_ed01]
signal BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2828_c7_006b]
signal t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2828_c7_006b]
signal t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2828_c7_006b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2828_c7_006b]
signal result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2828_c7_006b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2828_c7_006b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2828_c7_006b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2831_c11_697b]
signal BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2831_c7_5599]
signal t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2831_c7_5599]
signal t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2831_c7_5599]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2831_c7_5599]
signal result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2831_c7_5599]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2831_c7_5599]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2831_c7_5599]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2833_c30_f5a6]
signal sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2838_c11_0f3c]
signal BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2838_c7_72cc]
signal t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2838_c7_72cc]
signal result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2838_c7_72cc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2838_c7_72cc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2838_c7_72cc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2844_c11_d3dd]
signal BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2844_c7_205b]
signal result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2844_c7_205b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2844_c7_205b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2848_c11_0733]
signal BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2848_c7_1705]
signal result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2848_c7_1705]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2848_c7_1705]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e
BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_left,
BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_right,
BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec
t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec
t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec
result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec
result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec
result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec
result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec
result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec
result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec
result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01
BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_left,
BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_right,
BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2828_c7_006b
t16_low_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2828_c7_006b
t16_high_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b
result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b
result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b
result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b
BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_left,
BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_right,
BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2831_c7_5599
t16_low_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2831_c7_5599
t16_high_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599
result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599
result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599
result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599
result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6
sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_ins,
sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_x,
sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_y,
sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c
BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_left,
BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_right,
BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc
t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_cond,
t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue,
t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse,
t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc
result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc
result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd
BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_left,
BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_right,
BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b
result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b
result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733
BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_left,
BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_right,
BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705
result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_cond,
result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705
result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output,
 t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output,
 t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output,
 t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output,
 sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output,
 t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2820_c3_e84b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2825_c3_0a7b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2829_c3_56bc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2835_c3_0523 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2840_c3_8e59 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2841_c3_7530 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2845_c3_0024 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2849_c3_c49d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2848_c7_1705_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2848_l2815_l2828_DUPLICATE_851d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2838_l2828_DUPLICATE_f018_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2828_l2831_DUPLICATE_56d4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2854_l2811_DUPLICATE_ab84_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2829_c3_56bc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2829_c3_56bc;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2825_c3_0a7b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2825_c3_0a7b;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2835_c3_0523 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2835_c3_0523;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2840_c3_8e59 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2840_c3_8e59;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2849_c3_c49d := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2849_c3_c49d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2841_c3_7530 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2841_c3_7530;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2820_c3_e84b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2820_c3_e84b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2845_c3_0024 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2845_c3_0024;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2815_c6_813e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2828_c11_ed01] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_left;
     BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output := BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2838_c11_0f3c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output := result.is_stack_index_flipped;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output := result.is_vram_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2848_c7_1705] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2848_c7_1705_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2831_c11_697b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2833_c30_f5a6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_ins;
     sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_x;
     sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output := sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2848_l2815_l2828_DUPLICATE_851d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2848_l2815_l2828_DUPLICATE_851d_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2838_l2828_DUPLICATE_f018 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2838_l2828_DUPLICATE_f018_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2828_l2831_DUPLICATE_56d4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2828_l2831_DUPLICATE_56d4_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2848_c11_0733] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_left;
     BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output := BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2844_c11_d3dd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2815_c6_813e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2828_c11_ed01_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2831_c11_697b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2838_c11_0f3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2844_c11_d3dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2848_c11_0733_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2838_l2828_DUPLICATE_f018_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2838_l2828_DUPLICATE_f018_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2828_l2848_l2844_l2838_l2831_DUPLICATE_b3bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2828_l2831_DUPLICATE_56d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2828_l2831_DUPLICATE_56d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2848_l2815_l2828_DUPLICATE_851d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2848_l2815_l2828_DUPLICATE_851d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2848_l2815_l2828_DUPLICATE_851d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2815_c2_1cec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2848_c7_1705_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2833_c30_f5a6_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2838_c7_72cc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2848_c7_1705] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2838_c7_72cc] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_cond;
     t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output := t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2848_c7_1705] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output := result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2848_c7_1705] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2848_c7_1705_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2848_c7_1705_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2848_c7_1705_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2844_c7_205b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2844_c7_205b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2844_c7_205b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2844_c7_205b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2844_c7_205b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2844_c7_205b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2838_c7_72cc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2838_c7_72cc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2838_c7_72cc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2838_c7_72cc_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2831_c7_5599] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2831_c7_5599_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2828_c7_006b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2828_c7_006b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2815_c2_1cec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2854_l2811_DUPLICATE_ab84 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2854_l2811_DUPLICATE_ab84_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2815_c2_1cec_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2854_l2811_DUPLICATE_ab84_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2854_l2811_DUPLICATE_ab84_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
