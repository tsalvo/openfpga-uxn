-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 31
entity dup_0CLK_d4b33a56 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_d4b33a56;
architecture arch of dup_0CLK_d4b33a56 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2772_c6_795d]
signal BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2772_c2_b643]
signal t8_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2772_c2_b643]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2785_c11_f4f4]
signal BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2785_c7_279c]
signal t8_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2785_c7_279c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2785_c7_279c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2785_c7_279c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2785_c7_279c]
signal result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2785_c7_279c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2786_c30_46c9]
signal sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2788_c11_fdb6]
signal BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2788_c7_f6b9]
signal t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2788_c7_f6b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2788_c7_f6b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2788_c7_f6b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2788_c7_f6b9]
signal result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2788_c7_f6b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2794_c11_4232]
signal BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2794_c7_3e90]
signal result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2794_c7_3e90]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2794_c7_3e90]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d
BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_left,
BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_right,
BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output);

-- t8_MUX_uxn_opcodes_h_l2772_c2_b643
t8_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
t8_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
t8_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643
result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643
result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643
result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643
result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643
result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643
result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643
result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4
BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_left,
BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_right,
BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output);

-- t8_MUX_uxn_opcodes_h_l2785_c7_279c
t8_MUX_uxn_opcodes_h_l2785_c7_279c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2785_c7_279c_cond,
t8_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue,
t8_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse,
t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c
result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c
result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c
result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9
sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_ins,
sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_x,
sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_y,
sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6
BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_left,
BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_right,
BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output);

-- t8_MUX_uxn_opcodes_h_l2788_c7_f6b9
t8_MUX_uxn_opcodes_h_l2788_c7_f6b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond,
t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue,
t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse,
t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9
result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9
result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9
result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232
BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_left,
BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_right,
BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90
result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_cond,
result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90
result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output,
 t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output,
 t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output,
 t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2777_c3_41f1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2782_c3_f30a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2790_c3_faca : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2788_c7_f6b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2795_c3_b374 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2772_l2794_l2785_DUPLICATE_199e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_2a8a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2788_l2785_DUPLICATE_3999_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_ac10_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2800_l2768_DUPLICATE_4a98_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2777_c3_41f1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2777_c3_41f1;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2782_c3_f30a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2782_c3_f30a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2795_c3_b374 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2795_c3_b374;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2790_c3_faca := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2790_c3_faca;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_ac10 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_ac10_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2772_l2794_l2785_DUPLICATE_199e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2772_l2794_l2785_DUPLICATE_199e_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_2a8a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_2a8a_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2794_c11_4232] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_left;
     BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output := BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2788_l2785_DUPLICATE_3999 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2788_l2785_DUPLICATE_3999_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2772_c6_795d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2788_c11_fdb6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2785_c11_f4f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2772_c2_b643_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2772_c2_b643_return_output := result.is_pc_updated;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2788_c7_f6b9_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2786_c30_46c9] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_ins;
     sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_x;
     sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output := sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2772_c2_b643_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2772_c2_b643_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2772_c6_795d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2785_c11_f4f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2788_c11_fdb6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2794_c11_4232_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_ac10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_ac10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_ac10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2788_l2785_DUPLICATE_3999_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2788_l2785_DUPLICATE_3999_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_2a8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_2a8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2788_l2794_l2785_DUPLICATE_2a8a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2772_l2794_l2785_DUPLICATE_199e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2772_l2794_l2785_DUPLICATE_199e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2772_l2794_l2785_DUPLICATE_199e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2772_c2_b643_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2772_c2_b643_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2772_c2_b643_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2772_c2_b643_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2786_c30_46c9_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- t8_MUX[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond <= VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond;
     t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue;
     t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output := t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2794_c7_3e90] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2794_c7_3e90] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output := result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2794_c7_3e90] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2794_c7_3e90_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l2785_c7_279c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2785_c7_279c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_cond;
     t8_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue;
     t8_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output := t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2788_c7_f6b9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2785_c7_279c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2785_c7_279c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2788_c7_f6b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2785_c7_279c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2785_c7_279c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2785_c7_279c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     t8_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     t8_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2785_c7_279c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2772_c2_b643] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output;

     -- Submodule level 5
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2800_l2768_DUPLICATE_4a98 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2800_l2768_DUPLICATE_4a98_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2772_c2_b643_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2772_c2_b643_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2800_l2768_DUPLICATE_4a98_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2800_l2768_DUPLICATE_4a98_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
