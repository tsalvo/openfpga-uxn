-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity dup_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_66ba3dc0;
architecture arch of dup_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l3029_c6_5f75]
signal BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l3029_c1_c376]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3029_c2_7446]
signal t8_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3029_c2_7446]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3029_c2_7446]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3029_c2_7446]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3029_c2_7446]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3029_c2_7446]
signal result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3029_c2_7446]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l3030_c3_a95c[uxn_opcodes_h_l3030_c3_a95c]
signal printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3034_c11_3952]
signal BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3034_c7_2763]
signal t8_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3034_c7_2763]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3034_c7_2763]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3034_c7_2763]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3034_c7_2763]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3034_c7_2763]
signal result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3034_c7_2763]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3037_c11_794d]
signal BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3037_c7_6715]
signal t8_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3037_c7_6715]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3037_c7_6715]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3037_c7_6715]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3037_c7_6715]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3037_c7_6715]
signal result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3037_c7_6715]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l3040_c32_cfe4]
signal BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l3040_c32_9c4a]
signal BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l3040_c32_e956]
signal MUX_uxn_opcodes_h_l3040_c32_e956_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l3040_c32_e956_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3040_c32_e956_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3040_c32_e956_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3042_c11_eadf]
signal BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3042_c7_2431]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3042_c7_2431]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3042_c7_2431]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3042_c7_2431]
signal result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3042_c7_2431]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3048_c11_7022]
signal BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3048_c7_78a6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3048_c7_78a6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3048_c7_78a6]
signal result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3048_c7_78a6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3052_c11_0551]
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3052_c7_1b77]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3052_c7_1b77]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_53ff( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_value := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75
BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_left,
BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_right,
BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output);

-- t8_MUX_uxn_opcodes_h_l3029_c2_7446
t8_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
t8_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
t8_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446
result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446
result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446
result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446
result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446
result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

-- printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c
printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c : entity work.printf_uxn_opcodes_h_l3030_c3_a95c_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952
BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_left,
BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_right,
BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output);

-- t8_MUX_uxn_opcodes_h_l3034_c7_2763
t8_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
t8_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
t8_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763
result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763
result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763
result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763
result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763
result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d
BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_left,
BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_right,
BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output);

-- t8_MUX_uxn_opcodes_h_l3037_c7_6715
t8_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
t8_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
t8_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715
result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715
result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715
result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715
result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715
result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4
BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_left,
BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_right,
BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a
BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_left,
BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_right,
BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output);

-- MUX_uxn_opcodes_h_l3040_c32_e956
MUX_uxn_opcodes_h_l3040_c32_e956 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l3040_c32_e956_cond,
MUX_uxn_opcodes_h_l3040_c32_e956_iftrue,
MUX_uxn_opcodes_h_l3040_c32_e956_iffalse,
MUX_uxn_opcodes_h_l3040_c32_e956_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf
BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_left,
BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_right,
BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431
result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431
result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431
result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_cond,
result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431
result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022
BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_left,
BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_right,
BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6
result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6
result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_cond,
result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6
result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_left,
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_right,
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output,
 t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output,
 t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output,
 t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output,
 BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output,
 BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output,
 MUX_uxn_opcodes_h_l3040_c32_e956_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3031_c3_c8a7 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_3fa9 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3040_c32_e956_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3040_c32_e956_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3040_c32_e956_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3040_c32_e956_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3045_c3_495d : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_e65a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3037_l3029_l3034_DUPLICATE_a2ee_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3029_l3042_l3034_DUPLICATE_afae_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3037_l3048_DUPLICATE_4944_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l3057_l3025_DUPLICATE_7c2b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_e65a := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_e65a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3031_c3_c8a7 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3031_c3_c8a7;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_right := to_unsigned(128, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l3040_c32_e956_iffalse := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_MUX_uxn_opcodes_h_l3040_c32_e956_iftrue := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_right := to_unsigned(5, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_3fa9 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_3fa9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3045_c3_495d := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3045_c3_495d;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue := t8;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := t8;
     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3037_l3029_l3034_DUPLICATE_a2ee LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3037_l3029_l3034_DUPLICATE_a2ee_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l3048_c11_7022] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_left;
     BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output := BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3042_c11_eadf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_left;
     BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output := BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l3037_c11_794d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_left;
     BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output := BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3034_c11_3952] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_left;
     BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output := BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l3029_c6_5f75] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_left;
     BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output := BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3052_c11_0551] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_left;
     BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output := BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3037_l3048_DUPLICATE_4944 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3037_l3048_DUPLICATE_4944_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3029_l3042_l3034_DUPLICATE_afae LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3029_l3042_l3034_DUPLICATE_afae_return_output := result.is_sp_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l3040_c32_cfe4] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_left;
     BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output := BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_left := VAR_BIN_OP_AND_uxn_opcodes_h_l3040_c32_cfe4_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3029_c6_5f75_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3034_c11_3952_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3037_c11_794d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3042_c11_eadf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3048_c11_7022_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_0551_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3037_l3029_l3034_DUPLICATE_a2ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3037_l3029_l3034_DUPLICATE_a2ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3037_l3029_l3034_DUPLICATE_a2ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3037_l3034_l3052_l3048_l3042_DUPLICATE_4971_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3029_l3042_l3034_DUPLICATE_afae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3029_l3042_l3034_DUPLICATE_afae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3029_l3042_l3034_DUPLICATE_afae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3037_l3034_l3029_l3052_l3048_DUPLICATE_48ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3037_l3048_DUPLICATE_4944_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3037_l3048_DUPLICATE_4944_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3037_l3029_l3034_l3048_DUPLICATE_98ae_return_output;
     -- t8_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     t8_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     t8_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3048_c7_78a6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3048_c7_78a6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output := result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3052_c7_1b77] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3052_c7_1b77] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l3040_c32_9c4a] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_left;
     BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output := BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l3029_c1_c376] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3042_c7_2431] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l3040_c32_e956_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l3040_c32_9c4a_return_output;
     VAR_printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3029_c1_c376_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_1b77_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     -- printf_uxn_opcodes_h_l3030_c3_a95c[uxn_opcodes_h_l3030_c3_a95c] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l3030_c3_a95c_uxn_opcodes_h_l3030_c3_a95c_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3042_c7_2431] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3048_c7_78a6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3048_c7_78a6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;

     -- t8_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     t8_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     t8_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- MUX[uxn_opcodes_h_l3040_c32_e956] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l3040_c32_e956_cond <= VAR_MUX_uxn_opcodes_h_l3040_c32_e956_cond;
     MUX_uxn_opcodes_h_l3040_c32_e956_iftrue <= VAR_MUX_uxn_opcodes_h_l3040_c32_e956_iftrue;
     MUX_uxn_opcodes_h_l3040_c32_e956_iffalse <= VAR_MUX_uxn_opcodes_h_l3040_c32_e956_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l3040_c32_e956_return_output := MUX_uxn_opcodes_h_l3040_c32_e956_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3042_c7_2431] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output := result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue := VAR_MUX_uxn_opcodes_h_l3040_c32_e956_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3048_c7_78a6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l3042_c7_2431] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- t8_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     t8_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     t8_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3042_c7_2431] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3042_c7_2431_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3037_c7_6715] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3037_c7_6715_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3034_c7_2763] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3034_c7_2763_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3029_c2_7446] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l3057_l3025_DUPLICATE_7c2b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l3057_l3025_DUPLICATE_7c2b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_53ff(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3029_c2_7446_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3029_c2_7446_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l3057_l3025_DUPLICATE_7c2b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_53ff_uxn_opcodes_h_l3057_l3025_DUPLICATE_7c2b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
