-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity equ_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_85d5529e;
architecture arch of equ_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1114_c6_5582]
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1114_c1_6b10]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal n8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal t8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1114_c2_c02c]
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1115_c3_0e74[uxn_opcodes_h_l1115_c3_0e74]
signal printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1119_c11_a365]
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1119_c7_502f]
signal n8_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1119_c7_502f]
signal t8_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1119_c7_502f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1119_c7_502f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1119_c7_502f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1119_c7_502f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1119_c7_502f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1119_c7_502f]
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1122_c11_b4ca]
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1122_c7_559c]
signal n8_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1122_c7_559c]
signal t8_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1122_c7_559c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1122_c7_559c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1122_c7_559c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1122_c7_559c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1122_c7_559c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1122_c7_559c]
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1125_c11_016d]
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1125_c7_e7b9]
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1128_c30_97fa]
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1131_c21_c364]
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1131_c21_732d]
signal MUX_uxn_opcodes_h_l1131_c21_732d_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_732d_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_732d_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_732d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1133_c11_47c1]
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c7_d15b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c7_d15b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c7_d15b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_left,
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_right,
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output);

-- n8_MUX_uxn_opcodes_h_l1114_c2_c02c
n8_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- t8_MUX_uxn_opcodes_h_l1114_c2_c02c
t8_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

-- printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74
printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74 : entity work.printf_uxn_opcodes_h_l1115_c3_0e74_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_left,
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_right,
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output);

-- n8_MUX_uxn_opcodes_h_l1119_c7_502f
n8_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
n8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
n8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- t8_MUX_uxn_opcodes_h_l1119_c7_502f
t8_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
t8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
t8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_left,
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_right,
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output);

-- n8_MUX_uxn_opcodes_h_l1122_c7_559c
n8_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
n8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
n8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- t8_MUX_uxn_opcodes_h_l1122_c7_559c
t8_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
t8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
t8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_left,
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_right,
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output);

-- n8_MUX_uxn_opcodes_h_l1125_c7_e7b9
n8_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa
sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_ins,
sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_x,
sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_y,
sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_left,
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_right,
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output);

-- MUX_uxn_opcodes_h_l1131_c21_732d
MUX_uxn_opcodes_h_l1131_c21_732d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1131_c21_732d_cond,
MUX_uxn_opcodes_h_l1131_c21_732d_iftrue,
MUX_uxn_opcodes_h_l1131_c21_732d_iffalse,
MUX_uxn_opcodes_h_l1131_c21_732d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_left,
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_right,
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output,
 n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output,
 n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output,
 n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output,
 n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output,
 sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output,
 MUX_uxn_opcodes_h_l1131_c21_732d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_4df6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_9b9d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_4e7d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_732d_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_732d_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_732d_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_732d_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1122_l1125_DUPLICATE_e769_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1139_l1110_DUPLICATE_f021_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_y := resize(to_signed(-1, 2), 4);
     VAR_MUX_uxn_opcodes_h_l1131_c21_732d_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_4df6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_4df6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_4e7d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_4e7d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_9b9d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_9b9d;
     VAR_MUX_uxn_opcodes_h_l1131_c21_732d_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1114_c6_5582] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_left;
     BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output := BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1125_c11_016d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1131_c21_c364] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_left;
     BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output := BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1122_c11_b4ca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_left;
     BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output := BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1128_c30_97fa] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_ins;
     sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_x;
     sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output := sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1119_c11_a365] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_left;
     BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output := BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1122_l1125_DUPLICATE_e769 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1122_l1125_DUPLICATE_e769_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1133_c11_47c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_5582_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_a365_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_b4ca_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_016d_return_output;
     VAR_MUX_uxn_opcodes_h_l1131_c21_732d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_c364_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_47c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_44ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1133_l1122_l1125_l1119_DUPLICATE_fb98_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_c16f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1133_l1122_l1114_l1119_DUPLICATE_8760_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1122_l1125_DUPLICATE_e769_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1122_l1125_DUPLICATE_e769_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1122_l1114_l1125_l1119_DUPLICATE_6e13_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_97fa_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c7_d15b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output;

     -- MUX[uxn_opcodes_h_l1131_c21_732d] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1131_c21_732d_cond <= VAR_MUX_uxn_opcodes_h_l1131_c21_732d_cond;
     MUX_uxn_opcodes_h_l1131_c21_732d_iftrue <= VAR_MUX_uxn_opcodes_h_l1131_c21_732d_iftrue;
     MUX_uxn_opcodes_h_l1131_c21_732d_iffalse <= VAR_MUX_uxn_opcodes_h_l1131_c21_732d_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1131_c21_732d_return_output := MUX_uxn_opcodes_h_l1131_c21_732d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c7_d15b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c7_d15b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     t8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     t8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1114_c1_6b10] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue := VAR_MUX_uxn_opcodes_h_l1131_c21_732d_return_output;
     VAR_printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_6b10_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_d15b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     t8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     t8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- printf_uxn_opcodes_h_l1115_c3_0e74[uxn_opcodes_h_l1115_c3_0e74] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1115_c3_0e74_uxn_opcodes_h_l1115_c3_0e74_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     n8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     n8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1125_c7_e7b9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_e7b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     n8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     n8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1122_c7_559c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_559c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1119_c7_502f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_502f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1114_c2_c02c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1139_l1110_DUPLICATE_f021 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1139_l1110_DUPLICATE_f021_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_c02c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1139_l1110_DUPLICATE_f021_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1139_l1110_DUPLICATE_f021_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
