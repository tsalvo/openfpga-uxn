-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity ldz_0CLK_df07acae is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_df07acae;
architecture arch of ldz_0CLK_df07acae is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1557_c6_e874]
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1557_c1_7f0c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal t8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1557_c2_1e74]
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l1558_c3_0bf0[uxn_opcodes_h_l1558_c3_0bf0]
signal printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1562_c11_d34f]
signal BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1562_c7_8684]
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1562_c7_8684]
signal t8_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1562_c7_8684]
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1565_c11_7c47]
signal BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1565_c7_cfa0]
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(15 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1568_c32_1eb4]
signal BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1568_c32_ea60]
signal BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1568_c32_afc7]
signal MUX_uxn_opcodes_h_l1568_c32_afc7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1568_c32_afc7_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1568_c32_afc7_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1568_c32_afc7_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1571_c11_594c]
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(7 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1571_c7_5b28]
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1575_c11_c997]
signal BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1575_c7_416f]
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1575_c7_416f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1575_c7_416f]
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1575_c7_416f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1575_c7_416f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1581_c11_28fc]
signal BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1581_c7_3884]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1581_c7_3884]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b20( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_value := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.ram_addr := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_left,
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_right,
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74
tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- t8_MUX_uxn_opcodes_h_l1557_c2_1e74
t8_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

-- printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0
printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0 : entity work.printf_uxn_opcodes_h_l1558_c3_0bf0_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_left,
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_right,
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1562_c7_8684
tmp8_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- t8_MUX_uxn_opcodes_h_l1562_c7_8684
t8_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
t8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
t8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_left,
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_right,
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0
tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- t8_MUX_uxn_opcodes_h_l1565_c7_cfa0
t8_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4
BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_left,
BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_right,
BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60
BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_left,
BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_right,
BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output);

-- MUX_uxn_opcodes_h_l1568_c32_afc7
MUX_uxn_opcodes_h_l1568_c32_afc7 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1568_c32_afc7_cond,
MUX_uxn_opcodes_h_l1568_c32_afc7_iftrue,
MUX_uxn_opcodes_h_l1568_c32_afc7_iffalse,
MUX_uxn_opcodes_h_l1568_c32_afc7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_left,
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_right,
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28
tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_left,
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_right,
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1575_c7_416f
tmp8_MUX_uxn_opcodes_h_l1575_c7_416f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_cond,
tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue,
tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse,
tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_left,
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_right,
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output,
 tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output,
 MUX_uxn_opcodes_h_l1568_c32_afc7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output,
 tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iffalse : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_9e14 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1563_c3_6c9e : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_return_output : signed(7 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_732b_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1573_c21_3dff_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1578_c3_5130 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_da68_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1562_l1565_l1557_DUPLICATE_cdd8_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_60d4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1575_l1565_l1571_DUPLICATE_21e0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b20_uxn_opcodes_h_l1553_l1586_DUPLICATE_5007_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1578_c3_5130 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1578_c3_5130;
     VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_9e14 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_9e14;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_right := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1563_c3_6c9e := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1563_c3_6c9e;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_left := VAR_phase;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse := tmp8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1562_c11_d34f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1557_c6_e874] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_left;
     BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output := BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1575_c11_c997] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_left;
     BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output := BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1571_c11_594c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1573_c21_3dff] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1573_c21_3dff_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output := result.is_stack_write;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1562_l1565_l1557_DUPLICATE_cdd8 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1562_l1565_l1557_DUPLICATE_cdd8_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1581_c11_28fc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_left;
     BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output := BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_da68 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_da68_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1565_c11_7c47] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_left;
     BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output := BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1575_l1565_l1571_DUPLICATE_21e0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1575_l1565_l1571_DUPLICATE_21e0_return_output := result.stack_address_sp_offset;

     -- BIN_OP_AND[uxn_opcodes_h_l1568_c32_1eb4] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_left;
     BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output := BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1569_c21_732b] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_732b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_60d4 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_60d4_return_output := result.ram_addr;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_1eb4_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_e874_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_d34f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_7c47_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_594c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_c997_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_28fc_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_732b_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1573_c21_3dff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1562_l1565_l1557_DUPLICATE_cdd8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1562_l1565_l1557_DUPLICATE_cdd8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1562_l1565_l1557_DUPLICATE_cdd8_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_60d4_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_60d4_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_60d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1562_l1581_l1575_l1565_l1571_DUPLICATE_52e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_da68_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_da68_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1562_l1557_l1571_DUPLICATE_da68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1562_l1557_l1581_l1565_l1571_DUPLICATE_7063_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1575_l1565_l1571_DUPLICATE_21e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1575_l1565_l1571_DUPLICATE_21e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1575_l1565_l1571_DUPLICATE_21e0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1562_l1557_l1575_l1565_l1571_DUPLICATE_d659_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1575_c7_416f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1575_c7_416f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_cond;
     tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output := tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1581_c7_3884] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1575_c7_416f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1557_c1_7f0c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1581_c7_3884] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1568_c32_ea60] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_left;
     BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output := BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_ea60_return_output;
     VAR_printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1557_c1_7f0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_3884_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_3884_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1575_c7_416f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;

     -- MUX[uxn_opcodes_h_l1568_c32_afc7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1568_c32_afc7_cond <= VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_cond;
     MUX_uxn_opcodes_h_l1568_c32_afc7_iftrue <= VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_iftrue;
     MUX_uxn_opcodes_h_l1568_c32_afc7_iffalse <= VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_return_output := MUX_uxn_opcodes_h_l1568_c32_afc7_return_output;

     -- t8_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     t8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     t8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- printf_uxn_opcodes_h_l1558_c3_0bf0[uxn_opcodes_h_l1558_c3_0bf0] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1558_c3_0bf0_uxn_opcodes_h_l1558_c3_0bf0_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1575_c7_416f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue := VAR_MUX_uxn_opcodes_h_l1568_c32_afc7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_416f_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     -- result_ram_addr_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- t8_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1571_c7_5b28] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_5b28_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1565_c7_cfa0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_cfa0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1562_c7_8684] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_8684_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1557_c2_1e74] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b20_uxn_opcodes_h_l1553_l1586_DUPLICATE_5007 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b20_uxn_opcodes_h_l1553_l1586_DUPLICATE_5007_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b20(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output,
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_1e74_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b20_uxn_opcodes_h_l1553_l1586_DUPLICATE_5007_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b20_uxn_opcodes_h_l1553_l1586_DUPLICATE_5007_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
