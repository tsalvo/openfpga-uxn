-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc2_0CLK_180c5210 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_180c5210;
architecture arch of inc2_0CLK_180c5210 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_9a6b]
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1355_c2_9da5]
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_bb08]
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1368_c7_dfa9]
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_735e]
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1371_c7_06aa]
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_9b7c]
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output : unsigned(8 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1373_c30_8c28]
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_b7d0]
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_0a1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_0a1f]
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_0a1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_0a1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1378_c7_0a1f]
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_30c9]
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1379_c37_906e]
signal MUX_uxn_opcodes_h_l1379_c37_906e_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_906e_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_906e_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_906e_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_b174]
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_left,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_right,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5
t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5
t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_cond,
t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue,
t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse,
t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_left,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_right,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9
t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9
t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond,
t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue,
t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse,
t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_left,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_right,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa
t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa
t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_cond,
t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue,
t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse,
t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_left,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_right,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28
sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_ins,
sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_x,
sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_y,
sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_left,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_right,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f
t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond,
t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue,
t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse,
t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_left,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_right,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output);

-- MUX_uxn_opcodes_h_l1379_c37_906e
MUX_uxn_opcodes_h_l1379_c37_906e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1379_c37_906e_cond,
MUX_uxn_opcodes_h_l1379_c37_906e_iftrue,
MUX_uxn_opcodes_h_l1379_c37_906e_iffalse,
MUX_uxn_opcodes_h_l1379_c37_906e_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_left,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_right,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output,
 t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output,
 t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output,
 t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output,
 t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output,
 MUX_uxn_opcodes_h_l1379_c37_906e_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_2b2b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_3227 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_188a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_uxn_opcodes_h_l1372_c3_5625 : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_8622 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output : unsigned(8 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_7e1e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_0a1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_65da : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_uxn_opcodes_h_l1379_c3_4c69 : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_left : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_906e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_906e_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_906e_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_906e_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_1849_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4b16_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_41b3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_785d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1386_l1351_DUPLICATE_368a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_8622 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_8622;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_7e1e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_7e1e;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_2b2b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_2b2b;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_65da := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_65da;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l1379_c37_906e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_188a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_188a;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_3227 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_3227;
     VAR_MUX_uxn_opcodes_h_l1379_c37_906e_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_left := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_left := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse := t16_high;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_left := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := t16_low;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1378_c7_0a1f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_0a1f_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_785d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_785d_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_30c9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_41b3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_41b3_return_output := result.sp_relative_shift;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_9b7c] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_735e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_1849 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_1849_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4b16 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4b16_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_bb08] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_left;
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output := BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_b7d0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_9a6b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1373_c30_8c28] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_ins;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_x;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output := sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output := result.is_ram_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9a6b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_bb08_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_735e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_b7d0_return_output;
     VAR_MUX_uxn_opcodes_h_l1379_c37_906e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_30c9_return_output;
     VAR_t16_low_uxn_opcodes_h_l1372_c3_5625 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_9b7c_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_41b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_41b3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_785d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_785d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_785d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4b16_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4b16_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_1849_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_1849_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_1849_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_9da5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_0a1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8c28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_5625;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_5625;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_0a1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_0a1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_0a1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;

     -- MUX[uxn_opcodes_h_l1379_c37_906e] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1379_c37_906e_cond <= VAR_MUX_uxn_opcodes_h_l1379_c37_906e_cond;
     MUX_uxn_opcodes_h_l1379_c37_906e_iftrue <= VAR_MUX_uxn_opcodes_h_l1379_c37_906e_iftrue;
     MUX_uxn_opcodes_h_l1379_c37_906e_iffalse <= VAR_MUX_uxn_opcodes_h_l1379_c37_906e_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1379_c37_906e_return_output := MUX_uxn_opcodes_h_l1379_c37_906e_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_right := VAR_MUX_uxn_opcodes_h_l1379_c37_906e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_b174] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- Submodule level 3
     VAR_t16_high_uxn_opcodes_h_l1379_c3_4c69 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_b174_return_output, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_4c69;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_4c69;
     -- t16_low_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1378_c7_0a1f] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output := t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_0a1f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_0a1f_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_06aa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_06aa_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1368_c7_dfa9] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_cond;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output := t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_dfa9_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_9da5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;

     -- Submodule level 7
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1386_l1351_DUPLICATE_368a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1386_l1351_DUPLICATE_368a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_9da5_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1386_l1351_DUPLICATE_368a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1386_l1351_DUPLICATE_368a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
