-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_8d2aa467 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_8d2aa467;
architecture arch of sft_0CLK_8d2aa467 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2214_c6_f27b]
signal BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2214_c2_8271]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2214_c2_8271]
signal t8_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2214_c2_8271]
signal tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2214_c2_8271]
signal n8_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2227_c11_7bbc]
signal BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2227_c7_9810]
signal result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2227_c7_9810]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2227_c7_9810]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2227_c7_9810]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2227_c7_9810]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2227_c7_9810]
signal t8_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2227_c7_9810]
signal tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2227_c7_9810]
signal n8_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2230_c11_eceb]
signal BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2230_c7_e6f5]
signal n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2232_c30_057e]
signal sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2234_c11_ff28]
signal BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2234_c7_6d1c]
signal n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2237_c18_e113]
signal BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2237_c11_727f]
signal BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2237_c34_a50b]
signal CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2237_c11_b25a]
signal BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_243c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b
BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_left,
BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_right,
BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271
result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271
result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271
result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271
result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271
result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271
result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271
result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- t8_MUX_uxn_opcodes_h_l2214_c2_8271
t8_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
t8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
t8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2214_c2_8271
tmp8_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- n8_MUX_uxn_opcodes_h_l2214_c2_8271
n8_MUX_uxn_opcodes_h_l2214_c2_8271 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2214_c2_8271_cond,
n8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue,
n8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse,
n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc
BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_left,
BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_right,
BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810
result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810
result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810
result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810
result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- t8_MUX_uxn_opcodes_h_l2227_c7_9810
t8_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
t8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
t8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2227_c7_9810
tmp8_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- n8_MUX_uxn_opcodes_h_l2227_c7_9810
n8_MUX_uxn_opcodes_h_l2227_c7_9810 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2227_c7_9810_cond,
n8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue,
n8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse,
n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb
BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_left,
BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_right,
BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5
result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- t8_MUX_uxn_opcodes_h_l2230_c7_e6f5
t8_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5
tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- n8_MUX_uxn_opcodes_h_l2230_c7_e6f5
n8_MUX_uxn_opcodes_h_l2230_c7_e6f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond,
n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue,
n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse,
n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2232_c30_057e
sp_relative_shift_uxn_opcodes_h_l2232_c30_057e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_ins,
sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_x,
sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_y,
sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28
BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_left,
BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_right,
BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c
result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c
result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c
result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c
tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- n8_MUX_uxn_opcodes_h_l2234_c7_6d1c
n8_MUX_uxn_opcodes_h_l2234_c7_6d1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond,
n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue,
n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse,
n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113
BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_left,
BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_right,
BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f
BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_41db8d51 port map (
BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_left,
BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_right,
BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b
CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_x,
CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a
BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_ad8922d4 port map (
BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_left,
BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_right,
BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output,
 sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output,
 CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2224_c3_0a1f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2219_c3_8115 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2228_c3_bc6d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2239_c3_6d5b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2236_c3_606e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_eb4b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2227_l2234_DUPLICATE_1e49_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_7733_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2230_l2234_DUPLICATE_f244_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2210_l2244_DUPLICATE_e1c3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2239_c3_6d5b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2239_c3_6d5b;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2236_c3_606e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2236_c3_606e;
     VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2219_c3_8115 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2219_c3_8115;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2228_c3_bc6d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2228_c3_bc6d;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_right := to_unsigned(15, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2224_c3_0a1f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2224_c3_0a1f;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := tmp8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2230_l2234_DUPLICATE_f244 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2230_l2234_DUPLICATE_f244_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_eb4b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_eb4b_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2214_c2_8271_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2214_c6_f27b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;

     -- CONST_SR_4[uxn_opcodes_h_l2237_c34_a50b] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output := CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2214_c2_8271_return_output := result.is_ram_write;

     -- BIN_OP_AND[uxn_opcodes_h_l2237_c18_e113] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_left;
     BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output := BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_7733 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_7733_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2227_l2234_DUPLICATE_1e49 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2227_l2234_DUPLICATE_1e49_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2230_c11_eceb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2232_c30_057e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_ins;
     sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_x;
     sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output := sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2214_c2_8271_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2227_c11_7bbc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2234_c11_ff28] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_left;
     BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output := BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2214_c2_8271_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2237_c18_e113_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2214_c6_f27b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2227_c11_7bbc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c11_eceb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2234_c11_ff28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2227_l2234_DUPLICATE_1e49_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2227_l2234_DUPLICATE_1e49_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_7733_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_7733_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_7733_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_eb4b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_eb4b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2227_l2230_l2234_DUPLICATE_eb4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2230_l2234_DUPLICATE_f244_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2230_l2234_DUPLICATE_f244_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2227_l2230_l2214_l2234_DUPLICATE_4bcf_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_right := VAR_CONST_SR_4_uxn_opcodes_h_l2237_c34_a50b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2214_c2_8271_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2214_c2_8271_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2214_c2_8271_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2214_c2_8271_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2232_c30_057e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2237_c11_727f] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_left;
     BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output := BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- t8_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2237_c11_727f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     -- t8_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     t8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     t8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2237_c11_b25a] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_left;
     BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output := BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2237_c11_b25a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- t8_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     t8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     t8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- n8_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     n8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     n8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2234_c7_6d1c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2234_c7_6d1c_return_output;
     -- n8_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     n8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     n8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2230_c7_e6f5] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_cond;
     tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output := tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2230_c7_e6f5_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2227_c7_9810] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output := result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2227_c7_9810_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2214_c2_8271] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_cond;
     tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output := tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2214_c2_8271_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2210_l2244_DUPLICATE_e1c3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2210_l2244_DUPLICATE_e1c3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_243c(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2214_c2_8271_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2214_c2_8271_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2210_l2244_DUPLICATE_e1c3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2210_l2244_DUPLICATE_e1c3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
