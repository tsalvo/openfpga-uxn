-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity mul_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_6be78140;
architecture arch of mul_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1940_c6_4ee2]
signal BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal n8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1940_c2_f5de]
signal t8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1947_c11_181a]
signal BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal n8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1947_c7_8f64]
signal t8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1950_c11_51e5]
signal BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1950_c7_b573]
signal n8_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1950_c7_b573]
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1950_c7_b573]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1950_c7_b573]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1950_c7_b573]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1950_c7_b573]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1950_c7_b573]
signal t8_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1953_c11_5ed6]
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1953_c7_ba12]
signal n8_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1953_c7_ba12]
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1953_c7_ba12]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1953_c7_ba12]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1953_c7_ba12]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1953_c7_ba12]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1956_c30_0fff]
signal sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1959_c21_06cc]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1961_c11_0049]
signal BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1961_c7_470a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1961_c7_470a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1961_c7_470a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2
BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_left,
BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_right,
BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output);

-- n8_MUX_uxn_opcodes_h_l1940_c2_f5de
n8_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de
result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de
result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de
result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de
result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- t8_MUX_uxn_opcodes_h_l1940_c2_f5de
t8_MUX_uxn_opcodes_h_l1940_c2_f5de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond,
t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue,
t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse,
t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a
BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_left,
BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_right,
BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output);

-- n8_MUX_uxn_opcodes_h_l1947_c7_8f64
n8_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64
result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64
result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64
result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64
result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- t8_MUX_uxn_opcodes_h_l1947_c7_8f64
t8_MUX_uxn_opcodes_h_l1947_c7_8f64 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond,
t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue,
t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse,
t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_left,
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_right,
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output);

-- n8_MUX_uxn_opcodes_h_l1950_c7_b573
n8_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
n8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
n8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- t8_MUX_uxn_opcodes_h_l1950_c7_b573
t8_MUX_uxn_opcodes_h_l1950_c7_b573 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1950_c7_b573_cond,
t8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue,
t8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse,
t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_left,
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_right,
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output);

-- n8_MUX_uxn_opcodes_h_l1953_c7_ba12
n8_MUX_uxn_opcodes_h_l1953_c7_ba12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1953_c7_ba12_cond,
n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue,
n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse,
n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_cond,
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff
sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_ins,
sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_x,
sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_y,
sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_left,
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_right,
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output,
 n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output,
 n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output,
 n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output,
 n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output,
 sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1944_c3_6a94 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1948_c3_1259 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l1959_c3_90fe : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1958_c3_7a35 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1962_c3_cfcf : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1950_l1953_DUPLICATE_5b0a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1936_l1967_DUPLICATE_3909_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1962_c3_cfcf := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1962_c3_cfcf;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1958_c3_7a35 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1958_c3_7a35;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1948_c3_1259 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1948_c3_1259;
     VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1944_c3_6a94 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1944_c3_6a94;
     VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1950_c11_51e5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1950_l1953_DUPLICATE_5b0a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1950_l1953_DUPLICATE_5b0a_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1956_c30_0fff] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_ins;
     sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_x;
     sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output := sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1961_c11_0049] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_left;
     BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output := BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1947_c11_181a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1959_c21_06cc] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1940_c6_4ee2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1953_c11_5ed6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1940_c6_4ee2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1947_c11_181a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_51e5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_5ed6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_0049_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l1959_c3_90fe := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1959_c21_06cc_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_7373_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1950_l1953_l1947_l1961_DUPLICATE_fc41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1950_l1940_l1947_l1961_DUPLICATE_9def_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1950_l1953_DUPLICATE_5b0a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1950_l1953_DUPLICATE_5b0a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1950_l1940_l1953_l1947_DUPLICATE_5c92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1956_c30_0fff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue := VAR_result_u8_value_uxn_opcodes_h_l1959_c3_90fe;
     -- n8_MUX[uxn_opcodes_h_l1953_c7_ba12] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1953_c7_ba12_cond <= VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_cond;
     n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue;
     n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output := n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;

     -- t8_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     t8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     t8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1961_c7_470a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1953_c7_ba12] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output := result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1961_c7_470a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1953_c7_ba12] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1961_c7_470a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_470a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_470a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_470a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1953_c7_ba12] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;

     -- n8_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     n8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     n8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- t8_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1953_c7_ba12] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1953_c7_ba12] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_ba12_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1950_c7_b573] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;

     -- t8_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- n8_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_b573_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- n8_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1947_c7_8f64] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1947_c7_8f64_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1940_c2_f5de] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1936_l1967_DUPLICATE_3909 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1936_l1967_DUPLICATE_3909_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1940_c2_f5de_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1936_l1967_DUPLICATE_3909_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1936_l1967_DUPLICATE_3909_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
