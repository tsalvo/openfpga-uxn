-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2230_c6_c08a]
signal BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2230_c2_6a6d]
signal t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2243_c11_3799]
signal BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal n8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2243_c7_d39d]
signal t8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2246_c11_ae20]
signal BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal n8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2246_c7_cb38]
signal t8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2248_c30_d00a]
signal sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2250_c11_8e7e]
signal BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal n8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2250_c7_1b07]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2253_c18_7e81]
signal BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2253_c11_dc4c]
signal BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2253_c34_dce8]
signal CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2253_c11_ccbe]
signal BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a
BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_left,
BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_right,
BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d
tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- n8_MUX_uxn_opcodes_h_l2230_c2_6a6d
n8_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d
result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- t8_MUX_uxn_opcodes_h_l2230_c2_6a6d
t8_MUX_uxn_opcodes_h_l2230_c2_6a6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond,
t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue,
t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse,
t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799
BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_left,
BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_right,
BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d
tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- n8_MUX_uxn_opcodes_h_l2243_c7_d39d
n8_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d
result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d
result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d
result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- t8_MUX_uxn_opcodes_h_l2243_c7_d39d
t8_MUX_uxn_opcodes_h_l2243_c7_d39d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond,
t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue,
t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse,
t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20
BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_left,
BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_right,
BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38
tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- n8_MUX_uxn_opcodes_h_l2246_c7_cb38
n8_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38
result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38
result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38
result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38
result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- t8_MUX_uxn_opcodes_h_l2246_c7_cb38
t8_MUX_uxn_opcodes_h_l2246_c7_cb38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond,
t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue,
t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse,
t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a
sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_ins,
sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_x,
sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_y,
sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e
BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_left,
BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_right,
BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07
tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- n8_MUX_uxn_opcodes_h_l2250_c7_1b07
n8_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07
result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07
result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07
result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07
result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81
BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_left,
BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_right,
BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c
BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_left,
BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_right,
BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8
CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_x,
CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe
BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_left,
BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_right,
BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output,
 tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output,
 tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output,
 tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output,
 sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output,
 tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output,
 CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_37e2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2240_c3_9f63 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2244_c3_3186 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2252_c3_3207 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2255_c3_d6ec : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_0851_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2250_l2243_DUPLICATE_31e3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_4c44_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2246_l2250_DUPLICATE_f4bb_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2260_l2226_DUPLICATE_e8ff_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_right := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_right := to_unsigned(15, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2252_c3_3207 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2252_c3_3207;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2255_c3_d6ec := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2255_c3_d6ec;
     VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_37e2 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_37e2;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2240_c3_9f63 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2240_c3_9f63;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2244_c3_3186 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2244_c3_3186;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2246_c11_ae20] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_left;
     BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output := BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_0851 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_0851_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2246_l2250_DUPLICATE_f4bb LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2246_l2250_DUPLICATE_f4bb_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2250_c11_8e7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;

     -- CONST_SR_4[uxn_opcodes_h_l2253_c34_dce8] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output := CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_4c44 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_4c44_return_output := result.is_stack_write;

     -- BIN_OP_AND[uxn_opcodes_h_l2253_c18_7e81] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_left;
     BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output := BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2248_c30_d00a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_ins;
     sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_x;
     sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output := sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2243_c11_3799] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_left;
     BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output := BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2250_l2243_DUPLICATE_31e3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2250_l2243_DUPLICATE_31e3_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2230_c6_c08a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2253_c18_7e81_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2230_c6_c08a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2243_c11_3799_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2246_c11_ae20_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2250_c11_8e7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2250_l2243_DUPLICATE_31e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2250_l2243_DUPLICATE_31e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_0851_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_0851_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_0851_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_4c44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_4c44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2246_l2250_l2243_DUPLICATE_4c44_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2246_l2250_DUPLICATE_f4bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2246_l2250_DUPLICATE_f4bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2246_l2230_l2250_l2243_DUPLICATE_1499_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_right := VAR_CONST_SR_4_uxn_opcodes_h_l2253_c34_dce8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2248_c30_d00a_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- t8_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- n8_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2253_c11_dc4c] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_left;
     BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output := BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2253_c11_dc4c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     -- BIN_OP_SL[uxn_opcodes_h_l2253_c11_ccbe] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_left;
     BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output := BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- t8_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2253_c11_ccbe_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2250_c7_1b07] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_cond;
     tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output := tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2250_c7_1b07_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2246_c7_cb38] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_cond;
     tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output := tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2246_c7_cb38_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2243_c7_d39d] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_cond;
     tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output := tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2243_c7_d39d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2230_c2_6a6d] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_cond;
     tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output := tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2260_l2226_DUPLICATE_e8ff LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2260_l2226_DUPLICATE_e8ff_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2230_c2_6a6d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2260_l2226_DUPLICATE_e8ff_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2260_l2226_DUPLICATE_e8ff_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
