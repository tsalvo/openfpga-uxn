-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2175_c6_b1ee]
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2175_c2_2f00]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_2463]
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_e8b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2191_c11_04cb]
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2191_c7_9180]
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2191_c7_9180]
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2191_c7_9180]
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2191_c7_9180]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2191_c7_9180]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2191_c7_9180]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2191_c7_9180]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2193_c30_56d6]
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_879a]
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2198_c7_311b]
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_311b]
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_311b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_311b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_311b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_243c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_left,
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_right,
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00
t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00
t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_left,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_right,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3
t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3
t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_left,
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_right,
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2191_c7_9180
t16_low_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2191_c7_9180
t16_high_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6
sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_ins,
sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_x,
sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_y,
sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_left,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_right,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2198_c7_311b
t16_low_MUX_uxn_opcodes_h_l2198_c7_311b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_cond,
t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue,
t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse,
t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output,
 t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output,
 t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output,
 t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output,
 sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output,
 t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_ffd1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_367c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_636e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_3311 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_b65c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_cc0f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_311b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_1fed_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_4b02_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_8f43_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_8ea0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2206_l2171_DUPLICATE_8956_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_3311 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_3311;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_y := resize(to_signed(-2, 3), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_367c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_367c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_b65c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_b65c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_ffd1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_ffd1;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_cc0f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_cc0f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_636e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_636e;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse := t16_low;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2198_c7_311b] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_311b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_2463] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_left;
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output := BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_4b02 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_4b02_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2175_c6_b1ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_879a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_1fed LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_1fed_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_8ea0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_8ea0_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_8f43 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_8f43_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2191_c11_04cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l2193_c30_56d6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_ins;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_x;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output := sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_b1ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_2463_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_04cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_879a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_8f43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_8f43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_8ea0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_8ea0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_8ea0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_4b02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_4b02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_1fed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_1fed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2175_l2198_l2188_DUPLICATE_1fed_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_2f00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_311b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_56d6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_311b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_311b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2198_c7_311b] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_cond;
     t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output := t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_311b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_311b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_311b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2191_c7_9180] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output := result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_9180_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_e8b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_e8b3_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2175_c2_2f00] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_cond;
     t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output := t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2206_l2171_DUPLICATE_8956 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2206_l2171_DUPLICATE_8956_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_243c(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_2f00_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2206_l2171_DUPLICATE_8956_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2206_l2171_DUPLICATE_8956_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
