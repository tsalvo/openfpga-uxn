-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity dup_0CLK_5176672b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_5176672b;
architecture arch of dup_0CLK_5176672b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2448_c6_b56d]
signal BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2448_c2_142e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2448_c2_142e]
signal t8_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2448_c2_142e]
signal tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2455_c11_cb35]
signal BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2455_c7_d4b6]
signal tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2457_c30_6ad6]
signal sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2459_c11_a19f]
signal BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal t8_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2459_c7_45e0]
signal tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2462_c3_bf78]
signal CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2463_c3_2bd8]
signal BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2470_c11_3219]
signal BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2470_c7_cf9f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2470_c7_cf9f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2470_c7_cf9f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d
BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_left,
BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_right,
BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e
result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e
result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e
result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- t8_MUX_uxn_opcodes_h_l2448_c2_142e
t8_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
t8_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
t8_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2448_c2_142e
tmp16_MUX_uxn_opcodes_h_l2448_c2_142e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_cond,
tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue,
tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse,
tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_left,
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_right,
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- t8_MUX_uxn_opcodes_h_l2455_c7_d4b6
t8_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6
tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond,
tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue,
tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse,
tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6
sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_ins,
sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_x,
sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_y,
sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f
BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_left,
BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_right,
BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0
result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0
result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0
result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0
result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- t8_MUX_uxn_opcodes_h_l2459_c7_45e0
t8_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0
tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_cond,
tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue,
tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse,
tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78
CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_x,
CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8
BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_left,
BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_right,
BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_left,
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_right,
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f
result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output,
 sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output,
 CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2452_c3_9e6c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2467_c3_d24d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2459_l2448_DUPLICATE_5010_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2455_l2459_l2448_DUPLICATE_ee11_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_12ec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2448_DUPLICATE_d2f0_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_6ad2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2455_l2459_DUPLICATE_e5ae_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2470_l2455_l2459_DUPLICATE_5a24_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2461_l2463_DUPLICATE_9ba3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2476_l2443_DUPLICATE_d1e1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2452_c3_9e6c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2452_c3_9e6c;
     VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2467_c3_d24d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2467_c3_d24d;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_right := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := t8;
     VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := tmp16;
     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2461_l2463_DUPLICATE_9ba3 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2461_l2463_DUPLICATE_9ba3_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2459_c11_a19f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2457_c30_6ad6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_ins;
     sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_x;
     sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output := sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_12ec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_12ec_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2455_l2459_DUPLICATE_e5ae LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2455_l2459_DUPLICATE_e5ae_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2470_c11_3219] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_left;
     BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output := BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2459_l2448_DUPLICATE_5010 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2459_l2448_DUPLICATE_5010_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2448_DUPLICATE_d2f0 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2448_DUPLICATE_d2f0_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2470_l2455_l2459_DUPLICATE_5a24 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2470_l2455_l2459_DUPLICATE_5a24_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2448_c6_b56d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2455_l2459_l2448_DUPLICATE_ee11 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2455_l2459_l2448_DUPLICATE_ee11_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_6ad2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_6ad2_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2455_c11_cb35] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_left;
     BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output := BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c6_b56d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_cb35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2459_c11_a19f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_3219_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2461_l2463_DUPLICATE_9ba3_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2461_l2463_DUPLICATE_9ba3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2448_DUPLICATE_d2f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2448_DUPLICATE_d2f0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2455_l2459_l2448_DUPLICATE_ee11_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2455_l2459_l2448_DUPLICATE_ee11_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2455_l2459_l2448_DUPLICATE_ee11_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2470_l2455_l2459_DUPLICATE_5a24_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2470_l2455_l2459_DUPLICATE_5a24_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2470_l2455_l2459_DUPLICATE_5a24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2459_l2448_DUPLICATE_5010_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2459_l2448_DUPLICATE_5010_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_12ec_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_12ec_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_12ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_6ad2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_6ad2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2470_l2455_l2448_DUPLICATE_6ad2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2455_l2459_DUPLICATE_e5ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2455_l2459_DUPLICATE_e5ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2457_c30_6ad6_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2470_c7_cf9f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2462_c3_bf78] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output := CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output;

     -- t8_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2470_c7_cf9f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2470_c7_cf9f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output;

     -- Submodule level 2
     VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_left := VAR_CONST_SL_8_uxn_opcodes_h_l2462_c3_bf78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2470_c7_cf9f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2463_c3_2bd8] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_left;
     BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output := BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- Submodule level 3
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2463_c3_2bd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     t8_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     t8_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2459_c7_45e0] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_cond;
     tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output := tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2459_c7_45e0_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2455_c7_d4b6] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_cond;
     tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output := tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2455_c7_d4b6_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2448_c2_142e] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_cond;
     tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output := tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;

     -- Submodule level 6
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l2448_c2_142e_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2476_l2443_DUPLICATE_d1e1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2476_l2443_DUPLICATE_d1e1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c2_142e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2448_c2_142e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2476_l2443_DUPLICATE_d1e1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2476_l2443_DUPLICATE_d1e1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
