-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity sub2_0CLK_06b39b76 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end sub2_0CLK_06b39b76;
architecture arch of sub2_0CLK_06b39b76 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2248_c6_ba3c]
signal BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2248_c2_f8fa]
signal t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2256_c11_b159]
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2256_c7_9c9f]
signal t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2259_c11_9099]
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2259_c7_1f3b]
signal t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2262_c30_48f3]
signal sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2264_c11_5ea7]
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2264_c7_024b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2264_c7_024b]
signal result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2264_c7_024b]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2264_c7_024b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2264_c7_024b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2264_c7_024b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l2264_c7_024b]
signal n16_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2264_c7_024b]
signal tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(15 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2266_c11_3c57]
signal BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_left : unsigned(15 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_right : unsigned(15 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2272_c11_4e19]
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2272_c7_fb29]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2272_c7_fb29]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2272_c7_fb29]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c
BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_left,
BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_right,
BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa
result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- n16_MUX_uxn_opcodes_h_l2248_c2_f8fa
n16_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa
tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- t16_MUX_uxn_opcodes_h_l2248_c2_f8fa
t16_MUX_uxn_opcodes_h_l2248_c2_f8fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond,
t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue,
t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse,
t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_left,
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_right,
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- n16_MUX_uxn_opcodes_h_l2256_c7_9c9f
n16_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f
tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- t16_MUX_uxn_opcodes_h_l2256_c7_9c9f
t16_MUX_uxn_opcodes_h_l2256_c7_9c9f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond,
t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue,
t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse,
t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099
BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_left,
BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_right,
BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- n16_MUX_uxn_opcodes_h_l2259_c7_1f3b
n16_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b
tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- t16_MUX_uxn_opcodes_h_l2259_c7_1f3b
t16_MUX_uxn_opcodes_h_l2259_c7_1f3b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond,
t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue,
t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse,
t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3
sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_ins,
sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_x,
sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_y,
sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_left,
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_right,
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b
result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- n16_MUX_uxn_opcodes_h_l2264_c7_024b
n16_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
n16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
n16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2264_c7_024b
tmp16_MUX_uxn_opcodes_h_l2264_c7_024b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_cond,
tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue,
tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse,
tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57
BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57 : entity work.BIN_OP_MINUS_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_left,
BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_right,
BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_left,
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_right,
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2253_c3_a311 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2257_c3_bf5c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2269_c3_9b39 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2256_l2248_l2264_DUPLICATE_181f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2259_l2248_DUPLICATE_a2d5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2259_l2264_DUPLICATE_213c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2278_l2244_DUPLICATE_0e57_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_right := to_unsigned(2, 2);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2257_c3_bf5c := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2257_c3_bf5c;
     VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2269_c3_9b39 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2269_c3_9b39;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2253_c3_a311 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2253_c3_a311;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_right := to_unsigned(4, 3);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := t16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := tmp16;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2264_c11_5ea7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2259_c11_9099] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_left;
     BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output := BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2256_c11_b159] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_left;
     BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output := BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2259_l2248_DUPLICATE_a2d5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2259_l2248_DUPLICATE_a2d5_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2256_l2248_l2264_DUPLICATE_181f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2256_l2248_l2264_DUPLICATE_181f_return_output := result.is_sp_shift;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2266_c11_3c57] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2248_c6_ba3c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2272_c11_4e19] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_left;
     BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output := BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2259_l2264_DUPLICATE_213c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2259_l2264_DUPLICATE_213c_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l2262_c30_48f3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_ins;
     sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_x;
     sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output := sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2248_c6_ba3c_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_b159_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c11_9099_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_5ea7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_4e19_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2266_c11_3c57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2259_l2248_DUPLICATE_a2d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2259_l2248_DUPLICATE_a2d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2259_l2248_DUPLICATE_a2d5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2256_l2259_l2248_l2264_DUPLICATE_54a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_1114_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2256_l2248_l2264_DUPLICATE_181f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2256_l2248_l2264_DUPLICATE_181f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2256_l2248_l2264_DUPLICATE_181f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2264_DUPLICATE_8ad4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2272_l2259_l2248_DUPLICATE_54c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2259_l2264_DUPLICATE_213c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2259_l2264_DUPLICATE_213c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2262_c30_48f3_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2272_c7_fb29] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2272_c7_fb29] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output;

     -- t16_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- n16_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     n16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     n16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2272_c7_fb29] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_fb29_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- t16_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- n16_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2264_c7_024b] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_024b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     -- t16_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- n16_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2259_c7_1f3b] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c7_1f3b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- n16_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2256_c7_9c9f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_9c9f_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2248_c2_f8fa] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2278_l2244_DUPLICATE_0e57 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2278_l2244_DUPLICATE_0e57_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2248_c2_f8fa_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2278_l2244_DUPLICATE_0e57_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2278_l2244_DUPLICATE_0e57_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
