-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity nip_0CLK_6481cb28 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip_0CLK_6481cb28;
architecture arch of nip_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2425_c6_2574]
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2425_c1_bc5f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2425_c2_7fa7]
signal t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2426_c3_a120[uxn_opcodes_h_l2426_c3_a120]
signal printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2431_c11_ab2b]
signal BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2431_c7_16f4]
signal t8_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2434_c11_2623]
signal BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2434_c7_dbfa]
signal t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2438_c32_5dd2]
signal BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2438_c32_a19a]
signal BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2438_c32_1fd9]
signal MUX_uxn_opcodes_h_l2438_c32_1fd9_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2438_c32_1fd9_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2438_c32_1fd9_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2440_c11_328b]
signal BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2440_c7_9f47]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2440_c7_9f47]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2440_c7_9f47]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2440_c7_9f47]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2440_c7_9f47]
signal result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2446_c11_d42d]
signal BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2446_c7_ef9d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2446_c7_ef9d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_1ade( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.is_stack_read := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.stack_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_left,
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_right,
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7
result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- t8_MUX_uxn_opcodes_h_l2425_c2_7fa7
t8_MUX_uxn_opcodes_h_l2425_c2_7fa7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond,
t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue,
t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse,
t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

-- printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120
printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120 : entity work.printf_uxn_opcodes_h_l2426_c3_a120_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b
BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_left,
BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_right,
BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4
result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4
result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4
result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4
result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4
result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- t8_MUX_uxn_opcodes_h_l2431_c7_16f4
t8_MUX_uxn_opcodes_h_l2431_c7_16f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2431_c7_16f4_cond,
t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue,
t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse,
t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_left,
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_right,
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa
result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- t8_MUX_uxn_opcodes_h_l2434_c7_dbfa
t8_MUX_uxn_opcodes_h_l2434_c7_dbfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond,
t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue,
t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse,
t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2
BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_left,
BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_right,
BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a
BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_left,
BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_right,
BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output);

-- MUX_uxn_opcodes_h_l2438_c32_1fd9
MUX_uxn_opcodes_h_l2438_c32_1fd9 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2438_c32_1fd9_cond,
MUX_uxn_opcodes_h_l2438_c32_1fd9_iftrue,
MUX_uxn_opcodes_h_l2438_c32_1fd9_iffalse,
MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_left,
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_right,
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47
result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47
result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_cond,
result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_left,
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_right,
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output,
 MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2428_c3_5c2f : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2432_c3_4fdc : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2443_c3_4a07 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2425_l2440_l2431_DUPLICATE_b652_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2431_l2434_DUPLICATE_f3e3_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2431_l2434_DUPLICATE_e4bc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2440_l2434_DUPLICATE_8ef8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l2451_l2421_DUPLICATE_8a12_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_right := to_unsigned(1, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2432_c3_4fdc := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2432_c3_4fdc;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2428_c3_5c2f := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2428_c3_5c2f;
     VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_right := to_unsigned(128, 8);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2443_c3_4a07 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2443_c3_4a07;
     VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_iffalse := resize(to_signed(-1, 2), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2425_c6_2574] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_left;
     BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output := BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2431_c11_ab2b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2440_l2434_DUPLICATE_8ef8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2440_l2434_DUPLICATE_8ef8_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2434_c11_2623] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_left;
     BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output := BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2425_l2440_l2431_DUPLICATE_b652 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2425_l2440_l2431_DUPLICATE_b652_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2431_l2434_DUPLICATE_e4bc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2431_l2434_DUPLICATE_e4bc_return_output := result.is_stack_read;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16_return_output := result.stack_value;

     -- BIN_OP_AND[uxn_opcodes_h_l2438_c32_5dd2] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_left;
     BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output := BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2446_c11_d42d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2440_c11_328b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2431_l2434_DUPLICATE_f3e3 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2431_l2434_DUPLICATE_f3e3_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2438_c32_5dd2_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_2574_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2431_c11_ab2b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_2623_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_328b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_d42d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2431_l2434_DUPLICATE_f3e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2431_l2434_DUPLICATE_f3e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2431_l2434_DUPLICATE_f3e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2431_l2446_l2434_DUPLICATE_90e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2425_l2440_l2431_DUPLICATE_b652_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2425_l2440_l2431_DUPLICATE_b652_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2425_l2440_l2431_DUPLICATE_b652_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2431_l2434_DUPLICATE_e4bc_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2431_l2434_DUPLICATE_e4bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2431_l2446_l2434_DUPLICATE_ea1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2440_l2434_DUPLICATE_8ef8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2440_l2434_DUPLICATE_8ef8_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2425_l2440_l2431_l2434_DUPLICATE_8b16_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l2440_c7_9f47] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output := result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2446_c7_ef9d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2446_c7_ef9d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2440_c7_9f47] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2440_c7_9f47] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;

     -- t8_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2425_c1_bc5f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2438_c32_a19a] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_left;
     BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output := BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2438_c32_a19a_return_output;
     VAR_printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2425_c1_bc5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_ef9d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2440_c7_9f47] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;

     -- printf_uxn_opcodes_h_l2426_c3_a120[uxn_opcodes_h_l2426_c3_a120] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2426_c3_a120_uxn_opcodes_h_l2426_c3_a120_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2440_c7_9f47] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- MUX[uxn_opcodes_h_l2438_c32_1fd9] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2438_c32_1fd9_cond <= VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_cond;
     MUX_uxn_opcodes_h_l2438_c32_1fd9_iftrue <= VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_iftrue;
     MUX_uxn_opcodes_h_l2438_c32_1fd9_iffalse <= VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output := MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue := VAR_MUX_uxn_opcodes_h_l2438_c32_1fd9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_9f47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     -- t8_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2434_c7_dbfa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2434_c7_dbfa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2431_c7_16f4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2431_c7_16f4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c2_7fa7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l2451_l2421_DUPLICATE_8a12 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l2451_l2421_DUPLICATE_8a12_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1ade(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2425_c2_7fa7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l2451_l2421_DUPLICATE_8a12_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l2451_l2421_DUPLICATE_8a12_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
