-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_226c8821;
architecture arch of gth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_b4a1]
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1809_c2_8a8e]
signal t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_0e33]
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_5482]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_5482]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_5482]
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_5482]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_5482]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1822_c7_5482]
signal n8_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1822_c7_5482]
signal t8_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_1933]
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_7280]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_7280]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_7280]
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_7280]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_7280]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1825_c7_7280]
signal n8_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1825_c7_7280]
signal t8_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_901e]
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_357e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_357e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_357e]
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_357e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_357e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1828_c7_357e]
signal n8_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1830_c30_5fb5]
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1833_c21_e930]
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1833_c21_f30b]
signal MUX_uxn_opcodes_h_l1833_c21_f30b_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_f30b_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_f30b_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_f30b_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_left,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_right,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- n8_MUX_uxn_opcodes_h_l1809_c2_8a8e
n8_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- t8_MUX_uxn_opcodes_h_l1809_c2_8a8e
t8_MUX_uxn_opcodes_h_l1809_c2_8a8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond,
t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue,
t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse,
t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_left,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_right,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- n8_MUX_uxn_opcodes_h_l1822_c7_5482
n8_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
n8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
n8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- t8_MUX_uxn_opcodes_h_l1822_c7_5482
t8_MUX_uxn_opcodes_h_l1822_c7_5482 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1822_c7_5482_cond,
t8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue,
t8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse,
t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_left,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_right,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- n8_MUX_uxn_opcodes_h_l1825_c7_7280
n8_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
n8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
n8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- t8_MUX_uxn_opcodes_h_l1825_c7_7280
t8_MUX_uxn_opcodes_h_l1825_c7_7280 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1825_c7_7280_cond,
t8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue,
t8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse,
t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_left,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_right,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output);

-- n8_MUX_uxn_opcodes_h_l1828_c7_357e
n8_MUX_uxn_opcodes_h_l1828_c7_357e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1828_c7_357e_cond,
n8_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue,
n8_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse,
n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5
sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_ins,
sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_x,
sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_y,
sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_left,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_right,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output);

-- MUX_uxn_opcodes_h_l1833_c21_f30b
MUX_uxn_opcodes_h_l1833_c21_f30b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1833_c21_f30b_cond,
MUX_uxn_opcodes_h_l1833_c21_f30b_iftrue,
MUX_uxn_opcodes_h_l1833_c21_f30b_iffalse,
MUX_uxn_opcodes_h_l1833_c21_f30b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output,
 n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output,
 sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output,
 MUX_uxn_opcodes_h_l1833_c21_f30b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_ee55 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_2560 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_8b7d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_9bd9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f4c7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f60a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_db5d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_cdaf_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1837_l1805_DUPLICATE_8ba4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_2560 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_2560;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_y := resize(to_signed(-1, 2), 4);
     VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_8b7d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_8b7d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_9bd9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_9bd9;
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_ee55 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_ee55;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := t8;
     -- BIN_OP_GT[uxn_opcodes_h_l1833_c21_e930] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_left;
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output := BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_b4a1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_0e33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_left;
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output := BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_1933] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_left;
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output := BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_901e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output := result.is_vram_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_cdaf LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_cdaf_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1830_c30_5fb5] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_ins;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_x;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output := sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_db5d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_db5d_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f4c7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f4c7_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f60a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f60a_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_b4a1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_0e33_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1933_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_901e_return_output;
     VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e930_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f4c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f4c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f4c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_db5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_db5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_db5d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f60a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f60a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_f60a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_cdaf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_cdaf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1825_l1828_l1822_DUPLICATE_6879_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_8a8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_5fb5_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_357e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     t8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     t8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_357e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1828_c7_357e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1828_c7_357e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_cond;
     n8_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue;
     n8_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output := n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_357e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_357e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- MUX[uxn_opcodes_h_l1833_c21_f30b] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1833_c21_f30b_cond <= VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_cond;
     MUX_uxn_opcodes_h_l1833_c21_f30b_iftrue <= VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_iftrue;
     MUX_uxn_opcodes_h_l1833_c21_f30b_iffalse <= VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_return_output := MUX_uxn_opcodes_h_l1833_c21_f30b_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue := VAR_MUX_uxn_opcodes_h_l1833_c21_f30b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- n8_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     n8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     n8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- t8_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     t8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     t8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_357e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_357e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     -- n8_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     n8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     n8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_7280] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output := result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;

     -- t8_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_7280_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_5482] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output := result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_5482_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_8a8e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1837_l1805_DUPLICATE_8ba4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1837_l1805_DUPLICATE_8ba4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8a8e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1837_l1805_DUPLICATE_8ba4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1837_l1805_DUPLICATE_8ba4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
