-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_226c8821;
architecture arch of gth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1832_c6_6249]
signal BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal n8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal t8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1832_c2_4f30]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1845_c11_8e8f]
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1845_c7_6368]
signal n8_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1845_c7_6368]
signal t8_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1845_c7_6368]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1845_c7_6368]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1845_c7_6368]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1845_c7_6368]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1845_c7_6368]
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1848_c11_ce21]
signal BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal n8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal t8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1848_c7_36ee]
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1851_c11_bb77]
signal BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1851_c7_7dd2]
signal n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1851_c7_7dd2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1851_c7_7dd2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1851_c7_7dd2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1851_c7_7dd2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1851_c7_7dd2]
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1853_c30_a47c]
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1856_c21_d882]
signal BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1856_c21_f994]
signal MUX_uxn_opcodes_h_l1856_c21_f994_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1856_c21_f994_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1856_c21_f994_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1856_c21_f994_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e848( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_left,
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_right,
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output);

-- n8_MUX_uxn_opcodes_h_l1832_c2_4f30
n8_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- t8_MUX_uxn_opcodes_h_l1832_c2_4f30
t8_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_left,
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_right,
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output);

-- n8_MUX_uxn_opcodes_h_l1845_c7_6368
n8_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
n8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
n8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- t8_MUX_uxn_opcodes_h_l1845_c7_6368
t8_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
t8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
t8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_cond,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_left,
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_right,
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output);

-- n8_MUX_uxn_opcodes_h_l1848_c7_36ee
n8_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- t8_MUX_uxn_opcodes_h_l1848_c7_36ee
t8_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_cond,
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_left,
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_right,
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output);

-- n8_MUX_uxn_opcodes_h_l1851_c7_7dd2
n8_MUX_uxn_opcodes_h_l1851_c7_7dd2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond,
n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue,
n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse,
n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c
sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_ins,
sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_x,
sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_y,
sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882
BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_left,
BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_right,
BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output);

-- MUX_uxn_opcodes_h_l1856_c21_f994
MUX_uxn_opcodes_h_l1856_c21_f994 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1856_c21_f994_cond,
MUX_uxn_opcodes_h_l1856_c21_f994_iftrue,
MUX_uxn_opcodes_h_l1856_c21_f994_iffalse,
MUX_uxn_opcodes_h_l1856_c21_f994_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output,
 n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output,
 n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output,
 n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output,
 n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output,
 MUX_uxn_opcodes_h_l1856_c21_f994_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1837_c3_87b1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1842_c3_8f1d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1846_c3_66cb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1855_c3_0cd3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_f994_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_f994_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_f994_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_f994_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_69da_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_105a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_a460_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1848_l1851_DUPLICATE_57d9_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1860_l1828_DUPLICATE_1cc7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1842_c3_8f1d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1842_c3_8f1d;
     VAR_MUX_uxn_opcodes_h_l1856_c21_f994_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1855_c3_0cd3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1855_c3_0cd3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1837_c3_87b1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1837_c3_87b1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1846_c3_66cb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1846_c3_66cb;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1856_c21_f994_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1845_c11_8e8f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1832_c6_6249] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_left;
     BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output := BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1848_c11_ce21] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_left;
     BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output := BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1851_c11_bb77] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_left;
     BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output := BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_105a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_105a_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1853_c30_a47c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_ins;
     sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_x;
     sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output := sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1856_c21_d882] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_left;
     BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output := BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_a460 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_a460_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_69da LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_69da_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1848_l1851_DUPLICATE_57d9 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1848_l1851_DUPLICATE_57d9_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_6249_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_8e8f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_ce21_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_bb77_return_output;
     VAR_MUX_uxn_opcodes_h_l1856_c21_f994_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_d882_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_105a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_105a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_105a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_a460_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_a460_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_a460_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_69da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_69da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1848_l1851_l1845_DUPLICATE_69da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1848_l1851_DUPLICATE_57d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1848_l1851_DUPLICATE_57d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1848_l1832_l1851_l1845_DUPLICATE_660c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1832_c2_4f30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_a47c_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1851_c7_7dd2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1851_c7_7dd2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1851_c7_7dd2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond;
     n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue;
     n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output := n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1851_c7_7dd2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;

     -- MUX[uxn_opcodes_h_l1856_c21_f994] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1856_c21_f994_cond <= VAR_MUX_uxn_opcodes_h_l1856_c21_f994_cond;
     MUX_uxn_opcodes_h_l1856_c21_f994_iftrue <= VAR_MUX_uxn_opcodes_h_l1856_c21_f994_iftrue;
     MUX_uxn_opcodes_h_l1856_c21_f994_iffalse <= VAR_MUX_uxn_opcodes_h_l1856_c21_f994_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1856_c21_f994_return_output := MUX_uxn_opcodes_h_l1856_c21_f994_return_output;

     -- t8_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1851_c7_7dd2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue := VAR_MUX_uxn_opcodes_h_l1856_c21_f994_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     -- n8_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1851_c7_7dd2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- t8_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     t8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     t8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_7dd2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- t8_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- n8_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     n8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     n8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1848_c7_36ee] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output := result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_36ee_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1845_c7_6368] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output := result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;

     -- n8_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_6368_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1832_c2_4f30] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output := result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1860_l1828_DUPLICATE_1cc7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1860_l1828_DUPLICATE_1cc7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e848(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_4f30_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1860_l1828_DUPLICATE_1cc7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1860_l1828_DUPLICATE_1cc7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
