-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ovr_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_6d7675a8;
architecture arch of ovr_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l288_c6_9a3e]
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_94a5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l288_c2_809f]
signal n8_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l288_c2_809f]
signal t8_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_809f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_809f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_809f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_809f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_809f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l288_c2_809f]
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l289_c3_987a[uxn_opcodes_h_l289_c3_987a]
signal printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l293_c11_42a9]
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal n8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal t8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l293_c7_7e5b]
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l296_c11_68b1]
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal n8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal t8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l296_c7_2b8e]
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l299_c11_c135]
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l299_c7_c31d]
signal n8_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_c31d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_c31d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_c31d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_c31d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_c31d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l299_c7_c31d]
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l302_c30_b48a]
signal sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l307_c11_d35e]
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_667e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_667e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_667e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_667e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l307_c7_667e]
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l312_c11_5f54]
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_f7b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_f7b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_f7b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l312_c7_f7b6]
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l316_c11_b20d]
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_8468]
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_8468]
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e
BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_left,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_right,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output);

-- n8_MUX_uxn_opcodes_h_l288_c2_809f
n8_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l288_c2_809f_cond,
n8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
n8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- t8_MUX_uxn_opcodes_h_l288_c2_809f
t8_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l288_c2_809f_cond,
t8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
t8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f
result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_cond,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

-- printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a
printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a : entity work.printf_uxn_opcodes_h_l289_c3_987a_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9
BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_left,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_right,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output);

-- n8_MUX_uxn_opcodes_h_l293_c7_7e5b
n8_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- t8_MUX_uxn_opcodes_h_l293_c7_7e5b
t8_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b
result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_cond,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1
BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_left,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_right,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output);

-- n8_MUX_uxn_opcodes_h_l296_c7_2b8e
n8_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- t8_MUX_uxn_opcodes_h_l296_c7_2b8e
t8_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e
result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_cond,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135
BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_left,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_right,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output);

-- n8_MUX_uxn_opcodes_h_l299_c7_c31d
n8_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
n8_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
n8_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d
result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_cond,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l302_c30_b48a
sp_relative_shift_uxn_opcodes_h_l302_c30_b48a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_ins,
sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_x,
sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_y,
sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e
BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_left,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_right,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e
result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_cond,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_left,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_right,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6
result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d
BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_left,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_right,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output,
 n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output,
 n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output,
 n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output,
 n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output,
 sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_18a0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_3bde : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_ecf2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_a1a1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_65c0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_9bd8_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l321_l284_DUPLICATE_f32e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_a1a1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_a1a1;
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_3bde := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_3bde;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_65c0 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_65c0;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_18a0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_18a0;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_ecf2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_ecf2;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l296_c11_68b1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_left;
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output := BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l312_c11_5f54] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_left;
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output := BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l299_c11_c135] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_left;
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output := BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l288_c6_9a3e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_left;
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output := BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l293_c11_42a9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_left;
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output := BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l302_c30_b48a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_ins;
     sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_x;
     sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output := sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l307_c11_d35e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_left;
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output := BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_9bd8 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_9bd8_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l316_c11_b20d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_left;
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output := BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_9a3e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_42a9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_68b1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_c135_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_d35e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5f54_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_b20d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_a5d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l316_l312_l307_l299_l296_DUPLICATE_7346_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_fb70_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l316_l312_l307_l296_DUPLICATE_615a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_9bd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_9bd8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l288_l293_l296_DUPLICATE_d708_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_b48a_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_94a5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_8468] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_667e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- t8_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_8468] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l312_c7_f7b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;

     -- n8_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     n8_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     n8_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_f7b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_94a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_8468_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_667e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_8468_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     -- printf_uxn_opcodes_h_l289_c3_987a[uxn_opcodes_h_l289_c3_987a] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l289_c3_987a_uxn_opcodes_h_l289_c3_987a_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l307_c7_667e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output := result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_f7b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_667e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_f7b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;

     -- t8_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_f7b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_667e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_667e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     -- t8_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     t8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     t8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output := t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_667e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_667e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output;

     -- n8_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_667e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_667e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l288_c2_809f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- n8_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     n8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     n8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output := n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_c31d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l288_c2_809f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_c31d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_2b8e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_2b8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output := result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_7e5b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_7e5b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_809f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l321_l284_DUPLICATE_f32e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l321_l284_DUPLICATE_f32e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_809f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_809f_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l321_l284_DUPLICATE_f32e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l321_l284_DUPLICATE_f32e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
