-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity jcn_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jcn_0CLK_85d5529e;
architecture arch of jcn_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l644_c6_3810]
signal BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l644_c1_088a]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l644_c2_b3da]
signal t8_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l644_c2_b3da]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l644_c2_b3da]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l644_c2_b3da]
signal result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l644_c2_b3da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l644_c2_b3da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l644_c2_b3da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l644_c2_b3da]
signal n8_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l645_c3_0946[uxn_opcodes_h_l645_c3_0946]
signal printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l649_c11_6ac3]
signal BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l649_c7_ce16]
signal t8_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l649_c7_ce16]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l649_c7_ce16]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l649_c7_ce16]
signal result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l649_c7_ce16]
signal result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l649_c7_ce16]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l649_c7_ce16]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l649_c7_ce16]
signal n8_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l652_c11_6f82]
signal BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l652_c7_296b]
signal t8_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l652_c7_296b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l652_c7_296b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l652_c7_296b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l652_c7_296b]
signal result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l652_c7_296b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l652_c7_296b]
signal n8_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l655_c11_a2d0]
signal BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l655_c7_c7e7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l655_c7_c7e7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l655_c7_c7e7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l655_c7_c7e7]
signal result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l655_c7_c7e7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l655_c7_c7e7]
signal n8_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l658_c30_d585]
signal sp_relative_shift_uxn_opcodes_h_l658_c30_d585_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l658_c30_d585_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l658_c30_d585_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l660_c22_bb31]
signal BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l660_c37_b8c2]
signal BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output : signed(17 downto 0);

-- MUX[uxn_opcodes_h_l660_c22_7346]
signal MUX_uxn_opcodes_h_l660_c22_7346_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l660_c22_7346_iftrue : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l660_c22_7346_iffalse : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l660_c22_7346_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l662_c11_7833]
signal BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l662_c7_c4cc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l662_c7_c4cc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l662_c7_c4cc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a132( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810
BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_left,
BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_right,
BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output);

-- t8_MUX_uxn_opcodes_h_l644_c2_b3da
t8_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
t8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
t8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da
result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da
result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da
result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da
result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da
result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- n8_MUX_uxn_opcodes_h_l644_c2_b3da
n8_MUX_uxn_opcodes_h_l644_c2_b3da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l644_c2_b3da_cond,
n8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue,
n8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse,
n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

-- printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946
printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946 : entity work.printf_uxn_opcodes_h_l645_c3_0946_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3
BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_left,
BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_right,
BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output);

-- t8_MUX_uxn_opcodes_h_l649_c7_ce16
t8_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
t8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
t8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16
result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16
result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16
result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16
result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16
result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- n8_MUX_uxn_opcodes_h_l649_c7_ce16
n8_MUX_uxn_opcodes_h_l649_c7_ce16 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l649_c7_ce16_cond,
n8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue,
n8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse,
n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82
BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_left,
BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_right,
BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output);

-- t8_MUX_uxn_opcodes_h_l652_c7_296b
t8_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l652_c7_296b_cond,
t8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
t8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b
result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b
result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_cond,
result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- n8_MUX_uxn_opcodes_h_l652_c7_296b
n8_MUX_uxn_opcodes_h_l652_c7_296b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l652_c7_296b_cond,
n8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue,
n8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse,
n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0
BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_left,
BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_right,
BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7
result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7
result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7
result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7
result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_cond,
result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7
result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output);

-- n8_MUX_uxn_opcodes_h_l655_c7_c7e7
n8_MUX_uxn_opcodes_h_l655_c7_c7e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l655_c7_c7e7_cond,
n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue,
n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse,
n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l658_c30_d585
sp_relative_shift_uxn_opcodes_h_l658_c30_d585 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l658_c30_d585_ins,
sp_relative_shift_uxn_opcodes_h_l658_c30_d585_x,
sp_relative_shift_uxn_opcodes_h_l658_c30_d585_y,
sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31
BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_left,
BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_right,
BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2
BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_left,
BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_right,
BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output);

-- MUX_uxn_opcodes_h_l660_c22_7346
MUX_uxn_opcodes_h_l660_c22_7346 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l660_c22_7346_cond,
MUX_uxn_opcodes_h_l660_c22_7346_iftrue,
MUX_uxn_opcodes_h_l660_c22_7346_iffalse,
MUX_uxn_opcodes_h_l660_c22_7346_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833
BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_left,
BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_right,
BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output,
 t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output,
 t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output,
 t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output,
 n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output,
 sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output,
 MUX_uxn_opcodes_h_l660_c22_7346_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l646_c3_a5f8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l650_c3_89ce : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l649_c7_ce16_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l660_c22_7346_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l660_c22_7346_iftrue : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l660_c22_7346_iffalse : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l660_c42_78ca_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output : signed(17 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l660_c22_7346_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a132_uxn_opcodes_h_l668_l640_DUPLICATE_bbcf_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l646_c3_a5f8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l646_c3_a5f8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l650_c3_89ce := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l650_c3_89ce;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse := n8;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_MUX_uxn_opcodes_h_l660_c22_7346_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l652_c11_6f82] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_left;
     BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output := BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l658_c30_d585] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l658_c30_d585_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_ins;
     sp_relative_shift_uxn_opcodes_h_l658_c30_d585_x <= VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_x;
     sp_relative_shift_uxn_opcodes_h_l658_c30_d585_y <= VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output := sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l660_c22_bb31] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_left;
     BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output := BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l649_c11_6ac3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_left;
     BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output := BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l644_c6_3810] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_left;
     BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output := BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l662_c11_7833] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_left;
     BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output := BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l655_c11_a2d0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_left;
     BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output := BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l660_c42_78ca] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l660_c42_78ca_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l649_c7_ce16_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l644_c6_3810_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l649_c11_6ac3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c11_6f82_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l655_c11_a2d0_return_output;
     VAR_MUX_uxn_opcodes_h_l660_c22_7346_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c22_bb31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_7833_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l660_c42_78ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_3cbc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l644_l655_l649_l652_DUPLICATE_eb08_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l655_l649_l662_l652_DUPLICATE_9c71_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_f8f5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l644_l649_l662_l652_DUPLICATE_9b50_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l658_c30_d585_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l660_c37_b8c2] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_left;
     BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output := BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l662_c7_c4cc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l662_c7_c4cc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l662_c7_c4cc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output;

     -- t8_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     t8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     t8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output := t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- n8_MUX[uxn_opcodes_h_l655_c7_c7e7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l655_c7_c7e7_cond <= VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_cond;
     n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue;
     n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output := n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l644_c1_088a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l655_c7_c7e7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l660_c22_7346_iffalse := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l660_c37_b8c2_return_output)),16);
     VAR_printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l644_c1_088a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_c4cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_t8_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- n8_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     n8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     n8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output := n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l655_c7_c7e7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;

     -- MUX[uxn_opcodes_h_l660_c22_7346] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l660_c22_7346_cond <= VAR_MUX_uxn_opcodes_h_l660_c22_7346_cond;
     MUX_uxn_opcodes_h_l660_c22_7346_iftrue <= VAR_MUX_uxn_opcodes_h_l660_c22_7346_iftrue;
     MUX_uxn_opcodes_h_l660_c22_7346_iffalse <= VAR_MUX_uxn_opcodes_h_l660_c22_7346_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l660_c22_7346_return_output := MUX_uxn_opcodes_h_l660_c22_7346_return_output;

     -- printf_uxn_opcodes_h_l645_c3_0946[uxn_opcodes_h_l645_c3_0946] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l645_c3_0946_uxn_opcodes_h_l645_c3_0946_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l655_c7_c7e7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l655_c7_c7e7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;

     -- t8_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     t8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     t8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- Submodule level 3
     VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue := VAR_MUX_uxn_opcodes_h_l660_c22_7346_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_n8_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_t8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     -- t8_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     t8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     t8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- n8_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     n8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     n8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l655_c7_c7e7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output := result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_n8_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l655_c7_c7e7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l652_c7_296b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output := result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- n8_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     n8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     n8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c7_296b_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l649_c7_ce16] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_cond;
     result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output := result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- Submodule level 6
     VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l649_c7_ce16_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l644_c2_b3da] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_cond;
     result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output := result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a132_uxn_opcodes_h_l668_l640_DUPLICATE_bbcf LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a132_uxn_opcodes_h_l668_l640_DUPLICATE_bbcf_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a132(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l644_c2_b3da_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l644_c2_b3da_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a132_uxn_opcodes_h_l668_l640_DUPLICATE_bbcf_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a132_uxn_opcodes_h_l668_l640_DUPLICATE_bbcf_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
