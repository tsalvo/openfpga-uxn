-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity ovr_0CLK_12d025fa is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_12d025fa;
architecture arch of ovr_0CLK_12d025fa is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l300_c6_39fc]
signal BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l300_c2_5349]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l300_c2_5349]
signal n8_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l308_c11_39ac]
signal BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l308_c7_8624]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l308_c7_8624]
signal n8_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l310_c30_9e5f]
signal sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l312_c11_2bf4]
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_1f41]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l312_c7_1f41]
signal n8_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l313_c18_df7f]
signal CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l319_c11_0ea5]
signal BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l319_c7_270f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l319_c7_270f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l319_c7_270f]
signal result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l319_c7_270f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l319_c7_270f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l324_c11_6db6]
signal BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l324_c7_849f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l324_c7_849f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_4982( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_sp_shift := ref_toks_7;
      base.is_stack_operation_16bit := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc
BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_left,
BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_right,
BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349
result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349
result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349
result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349
result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349
result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349
result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- n8_MUX_uxn_opcodes_h_l300_c2_5349
n8_MUX_uxn_opcodes_h_l300_c2_5349 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l300_c2_5349_cond,
n8_MUX_uxn_opcodes_h_l300_c2_5349_iftrue,
n8_MUX_uxn_opcodes_h_l300_c2_5349_iffalse,
n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac
BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_left,
BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_right,
BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624
result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624
result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624
result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624
result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- n8_MUX_uxn_opcodes_h_l308_c7_8624
n8_MUX_uxn_opcodes_h_l308_c7_8624 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l308_c7_8624_cond,
n8_MUX_uxn_opcodes_h_l308_c7_8624_iftrue,
n8_MUX_uxn_opcodes_h_l308_c7_8624_iffalse,
n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output);

-- sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f
sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_ins,
sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_x,
sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_y,
sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4
BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_left,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_right,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41
result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41
result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41
result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- n8_MUX_uxn_opcodes_h_l312_c7_1f41
n8_MUX_uxn_opcodes_h_l312_c7_1f41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l312_c7_1f41_cond,
n8_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue,
n8_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse,
n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output);

-- CONST_SR_8_uxn_opcodes_h_l313_c18_df7f
CONST_SR_8_uxn_opcodes_h_l313_c18_df7f : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_x,
CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5
BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_left,
BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_right,
BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f
result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f
result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_cond,
result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f
result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6
BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_left,
BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_right,
BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f
result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f
result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output,
 sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output,
 CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_b079 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l316_c3_93ac : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l313_c8_4ad4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l321_c3_2c09 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l312_l300_l308_DUPLICATE_fbb7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l300_l308_DUPLICATE_4670_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l312_l300_DUPLICATE_cba7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l319_l308_DUPLICATE_ffb3_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l312_l319_l308_DUPLICATE_29ad_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l329_l296_DUPLICATE_5975_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_b079 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_b079;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l321_c3_2c09 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l321_c3_2c09;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l316_c3_93ac := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l316_c3_93ac;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_left := VAR_phase;
     VAR_CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_x := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := VAR_previous_stack_read;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l312_l300_DUPLICATE_cba7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l312_l300_DUPLICATE_cba7_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l312_l300_l308_DUPLICATE_fbb7 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l312_l300_l308_DUPLICATE_fbb7_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l312_l319_l308_DUPLICATE_29ad LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l312_l319_l308_DUPLICATE_29ad_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_EQ[uxn_opcodes_h_l324_c11_6db6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_left;
     BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output := BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l300_l308_DUPLICATE_4670 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l300_l308_DUPLICATE_4670_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l308_c11_39ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l319_c11_0ea5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_left;
     BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output := BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l319_l308_DUPLICATE_ffb3 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l319_l308_DUPLICATE_ffb3_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704_return_output := result.u8_value;

     -- CONST_SR_8[uxn_opcodes_h_l313_c18_df7f] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_x <= VAR_CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output := CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l310_c30_9e5f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_ins;
     sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_x;
     sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output := sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l312_c11_2bf4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_left;
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output := BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l300_c6_39fc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_left;
     BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output := BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l300_c6_39fc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_39ac_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_2bf4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l319_c11_0ea5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l324_c11_6db6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l300_l308_DUPLICATE_4670_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l300_l308_DUPLICATE_4670_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l312_l300_l308_DUPLICATE_fbb7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l312_l300_l308_DUPLICATE_fbb7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l312_l300_l308_DUPLICATE_fbb7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l324_l312_l319_l308_DUPLICATE_4b84_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l312_l300_DUPLICATE_cba7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l312_l300_DUPLICATE_cba7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l312_l319_l308_DUPLICATE_29ad_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l312_l319_l308_DUPLICATE_29ad_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l312_l319_l308_DUPLICATE_29ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l324_l300_l319_l308_DUPLICATE_c06d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l319_l308_DUPLICATE_ffb3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l319_l308_DUPLICATE_ffb3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l312_l300_l319_l308_DUPLICATE_9704_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_9e5f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l319_c7_270f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l319_c7_270f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l319_c7_270f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output := result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l324_c7_849f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l313_c8_4ad4] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l313_c8_4ad4_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l313_c18_df7f_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l324_c7_849f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l313_c8_4ad4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l324_c7_849f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l319_c7_270f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l324_c7_849f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l319_c7_270f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l319_c7_270f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- n8_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     n8_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     n8_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l319_c7_270f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l319_c7_270f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_n8_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l319_c7_270f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l319_c7_270f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_1f41] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- n8_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     n8_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     n8_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output := n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_n8_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_1f41_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- n8_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     n8_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     n8_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output := n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l308_c7_8624] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l300_c2_5349_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_8624_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l300_c2_5349] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l329_l296_DUPLICATE_5975 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l329_l296_DUPLICATE_5975_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4982(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l300_c2_5349_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l300_c2_5349_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l329_l296_DUPLICATE_5975_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l329_l296_DUPLICATE_5975_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
