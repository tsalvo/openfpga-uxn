-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity sub_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_fedec265;
architecture arch of sub_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2620_c6_d233]
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal n8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal t8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2620_c2_1a36]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2625_c11_7ae6]
signal BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2625_c7_750e]
signal n8_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2625_c7_750e]
signal t8_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2625_c7_750e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2625_c7_750e]
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2625_c7_750e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2625_c7_750e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2625_c7_750e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2625_c7_750e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2628_c11_d218]
signal BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal n8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal t8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2628_c7_39dc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2632_c11_8fc8]
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2632_c7_af36]
signal n8_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2632_c7_af36]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2632_c7_af36]
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2632_c7_af36]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2632_c7_af36]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2632_c7_af36]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2632_c7_af36]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2635_c11_3b30]
signal BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal n8_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2635_c7_9d38]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2638_c30_6e19]
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2641_c21_c935]
signal BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2643_c11_65c9]
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2643_c7_a8c9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2643_c7_a8c9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2643_c7_a8c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_left,
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_right,
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output);

-- n8_MUX_uxn_opcodes_h_l2620_c2_1a36
n8_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- t8_MUX_uxn_opcodes_h_l2620_c2_1a36
t8_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_left,
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_right,
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output);

-- n8_MUX_uxn_opcodes_h_l2625_c7_750e
n8_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
n8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
n8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- t8_MUX_uxn_opcodes_h_l2625_c7_750e
t8_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
t8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
t8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_left,
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_right,
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output);

-- n8_MUX_uxn_opcodes_h_l2628_c7_39dc
n8_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- t8_MUX_uxn_opcodes_h_l2628_c7_39dc
t8_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_left,
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_right,
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output);

-- n8_MUX_uxn_opcodes_h_l2632_c7_af36
n8_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
n8_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
n8_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_left,
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_right,
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output);

-- n8_MUX_uxn_opcodes_h_l2635_c7_9d38
n8_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19
sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_ins,
sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_x,
sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_y,
sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935
BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_left,
BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_right,
BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_left,
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_right,
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output,
 n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output,
 n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output,
 n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output,
 n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output,
 n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output,
 sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_f289 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_187b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2630_c3_a9c9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_d032 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_932b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2635_c7_9d38_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2616_l2649_DUPLICATE_dcc8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_187b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_187b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2630_c3_a9c9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2630_c3_a9c9;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_f289 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_f289;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_932b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_932b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_d032 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_d032;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2628_c11_d218] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_left;
     BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output := BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2641_c21_c935] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2632_c11_8fc8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2638_c30_6e19] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_ins;
     sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_x;
     sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output := sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2625_c11_7ae6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2635_c11_3b30] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_left;
     BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output := BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2635_c7_9d38_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2620_c6_d233] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_left;
     BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output := BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2643_c11_65c9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_d233_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_7ae6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_d218_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_8fc8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_3b30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_65c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2641_c21_c935_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_e5a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2643_l2635_DUPLICATE_193c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_ccd3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2643_DUPLICATE_40a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2628_l2625_l2620_l2635_DUPLICATE_b2ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_6e19_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- t8_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- n8_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2643_c7_a8c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2643_c7_a8c9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2643_c7_a8c9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_a8c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- n8_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     n8_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     n8_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- t8_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     t8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     t8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2635_c7_9d38] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_9d38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- n8_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- t8_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2632_c7_af36] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_af36_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     n8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     n8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2628_c7_39dc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_39dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2625_c7_750e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_750e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2620_c2_1a36] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2616_l2649_DUPLICATE_dcc8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2616_l2649_DUPLICATE_dcc8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_1a36_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2616_l2649_DUPLICATE_dcc8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2616_l2649_DUPLICATE_dcc8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
