-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity ora_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_bacf6a1d;
architecture arch of ora_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l956_c6_70fd]
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_d199]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal t8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l956_c2_5ed7]
signal n8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l957_c3_384e[uxn_opcodes_h_l957_c3_384e]
signal printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l961_c11_7131]
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l961_c7_5e77]
signal t8_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_5e77]
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_5e77]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_5e77]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_5e77]
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_5e77]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l961_c7_5e77]
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l961_c7_5e77]
signal n8_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l964_c11_98fb]
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l964_c7_7021]
signal t8_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_7021]
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_7021]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_7021]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_7021]
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_7021]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l964_c7_7021]
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l964_c7_7021]
signal n8_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l967_c11_2c5f]
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_7de0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_7de0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_7de0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_7de0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_7de0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l967_c7_7de0]
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l967_c7_7de0]
signal n8_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l970_c30_7fba]
signal sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l973_c21_9a2b]
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l975_c11_1fc1]
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_4fb6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_4fb6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_4fb6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd
BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_left,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_right,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output);

-- t8_MUX_uxn_opcodes_h_l956_c2_5ed7
t8_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7
result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- n8_MUX_uxn_opcodes_h_l956_c2_5ed7
n8_MUX_uxn_opcodes_h_l956_c2_5ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond,
n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue,
n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse,
n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

-- printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e
printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e : entity work.printf_uxn_opcodes_h_l957_c3_384e_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131
BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_left,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_right,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output);

-- t8_MUX_uxn_opcodes_h_l961_c7_5e77
t8_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
t8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
t8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77
result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- n8_MUX_uxn_opcodes_h_l961_c7_5e77
n8_MUX_uxn_opcodes_h_l961_c7_5e77 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l961_c7_5e77_cond,
n8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue,
n8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse,
n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb
BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_left,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_right,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output);

-- t8_MUX_uxn_opcodes_h_l964_c7_7021
t8_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l964_c7_7021_cond,
t8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
t8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021
result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_cond,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- n8_MUX_uxn_opcodes_h_l964_c7_7021
n8_MUX_uxn_opcodes_h_l964_c7_7021 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l964_c7_7021_cond,
n8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue,
n8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse,
n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f
BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_left,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_right,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0
result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- n8_MUX_uxn_opcodes_h_l967_c7_7de0
n8_MUX_uxn_opcodes_h_l967_c7_7de0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l967_c7_7de0_cond,
n8_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue,
n8_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse,
n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l970_c30_7fba
sp_relative_shift_uxn_opcodes_h_l970_c30_7fba : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_ins,
sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_x,
sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_y,
sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b
BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_left,
BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_right,
BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1
BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_left,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_right,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output,
 t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output,
 t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output,
 t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output,
 sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output,
 BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_7df8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_4e9f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_a55d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_b333_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l952_l981_DUPLICATE_0474_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_7df8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_7df8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_4e9f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_4e9f;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_y := resize(to_signed(-1, 2), 4);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_a55d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_a55d;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l975_c11_1fc1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_left;
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output := BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_b333 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_b333_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l970_c30_7fba] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_ins;
     sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_x <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_x;
     sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_y <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output := sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l967_c11_2c5f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_left;
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output := BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d_return_output := result.sp_relative_shift;

     -- BIN_OP_OR[uxn_opcodes_h_l973_c21_9a2b] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_left;
     BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output := BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l956_c6_70fd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_left;
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output := BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l964_c11_98fb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_left;
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output := BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l961_c11_7131] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_left;
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output := BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_70fd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_7131_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_98fb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_2c5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_1fc1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_9a2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_847d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_a6eb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2e3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_2c91_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_b333_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_b333_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_ded5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_7fba_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_4fb6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_d199] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_4fb6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_4fb6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- n8_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     n8_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     n8_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- t8_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     t8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     t8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output := t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_d199_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_n8_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4fb6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_t8_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     -- printf_uxn_opcodes_h_l957_c3_384e[uxn_opcodes_h_l957_c3_384e] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l957_c3_384e_uxn_opcodes_h_l957_c3_384e_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- t8_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     t8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     t8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_7de0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;

     -- n8_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     n8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     n8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output := n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output := result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_n8_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_7de0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- t8_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- n8_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     n8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     n8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_7021] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_7021_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- n8_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_5e77] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_5e77_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_5ed7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l952_l981_DUPLICATE_0474 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l952_l981_DUPLICATE_0474_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_5ed7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l952_l981_DUPLICATE_0474_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l952_l981_DUPLICATE_0474_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
