-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity and_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_f62d646e;
architecture arch of and_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l952_c6_636d]
signal BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l952_c1_f9f2]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l952_c2_1af7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l952_c2_1af7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l952_c2_1af7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l952_c2_1af7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l952_c2_1af7]
signal result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l952_c2_1af7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l952_c2_1af7]
signal t8_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l952_c2_1af7]
signal n8_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l953_c3_4364[uxn_opcodes_h_l953_c3_4364]
signal printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l957_c11_689d]
signal BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l957_c7_3f57]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l957_c7_3f57]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l957_c7_3f57]
signal result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l957_c7_3f57]
signal result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l957_c7_3f57]
signal result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l957_c7_3f57]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l957_c7_3f57]
signal t8_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l957_c7_3f57]
signal n8_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l960_c11_ab80]
signal BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l960_c7_1262]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l960_c7_1262]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l960_c7_1262]
signal result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l960_c7_1262]
signal result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l960_c7_1262]
signal result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l960_c7_1262]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l960_c7_1262]
signal t8_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l960_c7_1262]
signal n8_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l964_c11_9d61]
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_71a0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_71a0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_71a0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_71a0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l964_c7_71a0]
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_71a0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l964_c7_71a0]
signal n8_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l967_c11_fa47]
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l967_c7_1fa5]
signal n8_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l970_c30_ed93]
signal sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l973_c21_3aad]
signal BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l975_c11_d8c3]
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_4788]
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_4788]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_4788]
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d
BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_left,
BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_right,
BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7
result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7
result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7
result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- t8_MUX_uxn_opcodes_h_l952_c2_1af7
t8_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
t8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
t8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- n8_MUX_uxn_opcodes_h_l952_c2_1af7
n8_MUX_uxn_opcodes_h_l952_c2_1af7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l952_c2_1af7_cond,
n8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue,
n8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse,
n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

-- printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364
printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364 : entity work.printf_uxn_opcodes_h_l953_c3_4364_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d
BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_left,
BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_right,
BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57
result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57
result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57
result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57
result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57
result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- t8_MUX_uxn_opcodes_h_l957_c7_3f57
t8_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
t8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
t8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- n8_MUX_uxn_opcodes_h_l957_c7_3f57
n8_MUX_uxn_opcodes_h_l957_c7_3f57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l957_c7_3f57_cond,
n8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue,
n8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse,
n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80
BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_left,
BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_right,
BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262
result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262
result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262
result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262
result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_cond,
result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262
result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- t8_MUX_uxn_opcodes_h_l960_c7_1262
t8_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l960_c7_1262_cond,
t8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
t8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- n8_MUX_uxn_opcodes_h_l960_c7_1262
n8_MUX_uxn_opcodes_h_l960_c7_1262 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l960_c7_1262_cond,
n8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue,
n8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse,
n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_left,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_right,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0
result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- n8_MUX_uxn_opcodes_h_l964_c7_71a0
n8_MUX_uxn_opcodes_h_l964_c7_71a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l964_c7_71a0_cond,
n8_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue,
n8_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse,
n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47
BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_left,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_right,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5
result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- n8_MUX_uxn_opcodes_h_l967_c7_1fa5
n8_MUX_uxn_opcodes_h_l967_c7_1fa5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l967_c7_1fa5_cond,
n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue,
n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse,
n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output);

-- sp_relative_shift_uxn_opcodes_h_l970_c30_ed93
sp_relative_shift_uxn_opcodes_h_l970_c30_ed93 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_ins,
sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_x,
sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_y,
sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad
BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_left,
BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_right,
BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_left,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_right,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output,
 sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output,
 BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l954_c3_7db8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_a7b2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_ece5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l965_c3_e6e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_37d7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_c7_1fa5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l948_l981_DUPLICATE_d440_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l965_c3_e6e5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l965_c3_e6e5;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_a7b2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_a7b2;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l954_c3_7db8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l954_c3_7db8;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_37d7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_37d7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_ece5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_ece5;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l967_c11_fa47] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_left;
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output := BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l973_c21_3aad] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_left;
     BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output := BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l975_c11_d8c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l952_c6_636d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_left;
     BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output := BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l957_c11_689d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_left;
     BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output := BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l964_c11_9d61] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_left;
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output := BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l970_c30_ed93] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_ins;
     sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_x <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_x;
     sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_y <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output := sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l960_c11_ab80] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_left;
     BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output := BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_c7_1fa5_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l973_c21_3aad_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c6_636d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l957_c11_689d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l960_c11_ab80_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9d61_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_fa47_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d8c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_33ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l967_l964_l960_l957_DUPLICATE_78f6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_3cb8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l952_l975_l964_l960_l957_DUPLICATE_8dac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l952_l967_l964_l960_l957_DUPLICATE_1d08_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_ed93_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l952_c1_f9f2] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_4788] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output;

     -- n8_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_4788] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_4788] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output;

     -- t8_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     t8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     t8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output := t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l952_c1_f9f2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_4788_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_4788_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_4788_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_t8_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- n8_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     n8_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     n8_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- t8_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     t8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     t8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- printf_uxn_opcodes_h_l953_c3_4364[uxn_opcodes_h_l953_c3_4364] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l953_c3_4364_uxn_opcodes_h_l953_c3_4364_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_1fa5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_n8_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_1fa5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output := result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- n8_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     n8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     n8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output := n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- t8_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     t8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     t8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_71a0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_n8_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_71a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l960_c7_1262] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output;

     -- n8_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     n8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     n8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l960_c7_1262_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- n8_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     n8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     n8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l957_c7_3f57] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l957_c7_3f57_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l952_c2_1af7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l948_l981_DUPLICATE_d440 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l948_l981_DUPLICATE_d440_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c2_1af7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c2_1af7_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l948_l981_DUPLICATE_d440_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l948_l981_DUPLICATE_d440_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
