-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity opc_ovr_phased_0CLK_60e6c3c2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_ovr_phased_0CLK_60e6c3c2;
architecture arch of opc_ovr_phased_0CLK_60e6c3c2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l340_c6_e07a]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l340_c1_966f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l343_c7_b0dd]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l340_c2_b15f]
signal t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l340_c2_b15f]
signal n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l340_c2_b15f]
signal result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l341_c12_fcf7]
signal set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l343_c11_f475]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l343_c1_c11a]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l346_c7_d915]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l343_c7_b0dd]
signal t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l343_c7_b0dd]
signal n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l343_c7_b0dd]
signal result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l344_c8_b472]
signal t_register_uxn_opcodes_phased_h_l344_c8_b472_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l346_c11_b178]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l346_c1_c6a0]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l349_c7_789d]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l346_c7_d915]
signal t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l346_c7_d915]
signal n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l346_c7_d915]
signal result_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l347_c8_2927]
signal n_register_uxn_opcodes_phased_h_l347_c8_2927_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l349_c11_9b45]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l349_c1_1c10]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l352_c7_2df6]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l349_c7_789d]
signal n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l349_c7_789d]
signal result_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l350_c8_1c5b]
signal n_register_uxn_opcodes_phased_h_l350_c8_1c5b_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l352_c11_de7e]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l352_c1_9e3b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l355_c7_986d]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l352_c7_2df6]
signal result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l353_c3_8c81]
signal set_uxn_opcodes_phased_h_l353_c3_8c81_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l353_c3_8c81_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l353_c3_8c81_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l353_c3_8c81_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l353_c3_8c81_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l353_c3_8c81_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l353_c3_8c81_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l355_c11_9c3f]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l355_c1_06d3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l358_c7_d34c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l355_c7_986d]
signal result_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_phased_h_l356_c3_adfd]
signal put_stack_uxn_opcodes_phased_h_l356_c3_adfd_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l356_c3_adfd_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l356_c3_adfd_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l356_c3_adfd_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l356_c3_adfd_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l358_c11_3a2b]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l358_c1_f6de]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l361_c7_6668]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l358_c7_d34c]
signal result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_phased_h_l359_c3_2fb0]
signal put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l361_c11_15a7]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l361_c1_8ca3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l361_c7_6668]
signal result_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_phased_h_l362_c3_9e5b]
signal put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l364_c11_c3d1]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_right : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l364_c7_af44]
signal result_MUX_uxn_opcodes_phased_h_l364_c7_af44_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a
BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f
t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond,
t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue,
t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse,
t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f
n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond,
n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue,
n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse,
n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output);

-- result_MUX_uxn_opcodes_phased_h_l340_c2_b15f
result_MUX_uxn_opcodes_phased_h_l340_c2_b15f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond,
result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue,
result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse,
result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_sp,
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_k,
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_mul,
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_add,
set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475
BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd
t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond,
t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue,
t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse,
t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd
n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond,
n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue,
n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse,
n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output);

-- result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd
result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond,
result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue,
result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse,
result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output);

-- t_register_uxn_opcodes_phased_h_l344_c8_b472
t_register_uxn_opcodes_phased_h_l344_c8_b472 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l344_c8_b472_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_index,
t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_ptr,
t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178
BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l346_c7_d915
t8_MUX_uxn_opcodes_phased_h_l346_c7_d915 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond,
t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue,
t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse,
t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l346_c7_d915
n8_MUX_uxn_opcodes_phased_h_l346_c7_d915 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond,
n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue,
n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse,
n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output);

-- result_MUX_uxn_opcodes_phased_h_l346_c7_d915
result_MUX_uxn_opcodes_phased_h_l346_c7_d915 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond,
result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue,
result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse,
result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output);

-- n_register_uxn_opcodes_phased_h_l347_c8_2927
n_register_uxn_opcodes_phased_h_l347_c8_2927 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l347_c8_2927_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_index,
n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_ptr,
n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45
BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l349_c7_789d
n8_MUX_uxn_opcodes_phased_h_l349_c7_789d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond,
n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue,
n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse,
n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output);

-- result_MUX_uxn_opcodes_phased_h_l349_c7_789d
result_MUX_uxn_opcodes_phased_h_l349_c7_789d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond,
result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue,
result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse,
result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output);

-- n_register_uxn_opcodes_phased_h_l350_c8_1c5b
n_register_uxn_opcodes_phased_h_l350_c8_1c5b : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l350_c8_1c5b_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_index,
n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_ptr,
n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e
BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output);

-- result_MUX_uxn_opcodes_phased_h_l352_c7_2df6
result_MUX_uxn_opcodes_phased_h_l352_c7_2df6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond,
result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue,
result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse,
result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output);

-- set_uxn_opcodes_phased_h_l353_c3_8c81
set_uxn_opcodes_phased_h_l353_c3_8c81 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l353_c3_8c81_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l353_c3_8c81_sp,
set_uxn_opcodes_phased_h_l353_c3_8c81_stack_index,
set_uxn_opcodes_phased_h_l353_c3_8c81_ins,
set_uxn_opcodes_phased_h_l353_c3_8c81_k,
set_uxn_opcodes_phased_h_l353_c3_8c81_mul,
set_uxn_opcodes_phased_h_l353_c3_8c81_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f
BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l355_c7_986d
result_MUX_uxn_opcodes_phased_h_l355_c7_986d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond,
result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue,
result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse,
result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output);

-- put_stack_uxn_opcodes_phased_h_l356_c3_adfd
put_stack_uxn_opcodes_phased_h_l356_c3_adfd : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l356_c3_adfd_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l356_c3_adfd_sp,
put_stack_uxn_opcodes_phased_h_l356_c3_adfd_stack_index,
put_stack_uxn_opcodes_phased_h_l356_c3_adfd_offset,
put_stack_uxn_opcodes_phased_h_l356_c3_adfd_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b
BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output);

-- result_MUX_uxn_opcodes_phased_h_l358_c7_d34c
result_MUX_uxn_opcodes_phased_h_l358_c7_d34c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond,
result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue,
result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse,
result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output);

-- put_stack_uxn_opcodes_phased_h_l359_c3_2fb0
put_stack_uxn_opcodes_phased_h_l359_c3_2fb0 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_sp,
put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_stack_index,
put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_offset,
put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7
BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output);

-- result_MUX_uxn_opcodes_phased_h_l361_c7_6668
result_MUX_uxn_opcodes_phased_h_l361_c7_6668 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond,
result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue,
result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse,
result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output);

-- put_stack_uxn_opcodes_phased_h_l362_c3_9e5b
put_stack_uxn_opcodes_phased_h_l362_c3_9e5b : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_sp,
put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_stack_index,
put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_offset,
put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1
BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output);

-- result_MUX_uxn_opcodes_phased_h_l364_c7_af44
result_MUX_uxn_opcodes_phased_h_l364_c7_af44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l364_c7_af44_cond,
result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iftrue,
result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iffalse,
result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output,
 t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output,
 n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output,
 result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output,
 set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output,
 t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output,
 n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output,
 result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output,
 t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output,
 t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output,
 n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output,
 result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output,
 n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output,
 n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output,
 result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output,
 n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output,
 result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output,
 result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output,
 result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output,
 result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output,
 result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_right := to_unsigned(7, 3);
     VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_offset := resize(to_unsigned(2, 2), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_mul := resize(to_unsigned(2, 2), 8);
     VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue := to_unsigned(0, 1);
     VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_offset := resize(to_unsigned(0, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_add := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_right := to_unsigned(2, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_right := to_unsigned(5, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_add := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_right := to_unsigned(3, 2);
     VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_offset := resize(to_unsigned(1, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_k := VAR_k;
     VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse := n8;
     VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_value := n8;
     VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_value := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_sp := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_sp := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_value := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l364_c11_c3d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l361_c11_15a7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l343_c11_f475] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l352_c11_de7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l340_c6_e07a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l358_c11_3a2b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l346_c11_b178] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l355_c11_9c3f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l349_c11_9b45] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l340_c6_e07a_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l343_c11_f475_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l346_c11_b178_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l349_c11_9b45_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l352_c11_de7e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l355_c11_9c3f_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l358_c11_3a2b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l361_c11_15a7_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l364_c11_c3d1_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l343_c7_b0dd] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l364_c7_af44] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l364_c7_af44_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_cond;
     result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iftrue;
     result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output := result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l340_c1_966f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l340_c1_966f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l364_c7_af44_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l346_c7_d915] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l343_c1_c11a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l361_c7_6668] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond;
     result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue;
     result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output := result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l341_c12_fcf7] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_sp;
     set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_k;
     set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_mul;
     set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output := set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l343_c1_c11a_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l341_c12_fcf7_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l349_c7_789d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;

     -- t_register[uxn_opcodes_phased_h_l344_c8_b472] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l344_c8_b472_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_index;
     t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output := t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l346_c1_c6a0] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l358_c7_d34c] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond;
     result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue;
     result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output := result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l346_c1_c6a0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue := VAR_t_register_uxn_opcodes_phased_h_l344_c8_b472_return_output;
     -- n_register[uxn_opcodes_phased_h_l347_c8_2927] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l347_c8_2927_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_index;
     n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output := n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l349_c1_1c10] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l352_c7_2df6] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l355_c7_986d] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond;
     result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue;
     result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output := result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l349_c1_1c10_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue := VAR_n_register_uxn_opcodes_phased_h_l347_c8_2927_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l355_c7_986d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output;

     -- n_register[uxn_opcodes_phased_h_l350_c8_1c5b] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l350_c8_1c5b_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_index;
     n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output := n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l352_c1_9e3b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l346_c7_d915] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond;
     t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output := t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l352_c7_2df6] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_cond;
     result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iftrue;
     result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output := result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output;

     -- Submodule level 6
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c7_986d_return_output;
     VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l352_c1_9e3b_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue := VAR_n_register_uxn_opcodes_phased_h_l350_c8_1c5b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l352_c7_2df6_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;
     -- set[uxn_opcodes_phased_h_l353_c3_8c81] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l353_c3_8c81_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l353_c3_8c81_sp <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_sp;
     set_uxn_opcodes_phased_h_l353_c3_8c81_stack_index <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_stack_index;
     set_uxn_opcodes_phased_h_l353_c3_8c81_ins <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_ins;
     set_uxn_opcodes_phased_h_l353_c3_8c81_k <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_k;
     set_uxn_opcodes_phased_h_l353_c3_8c81_mul <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_mul;
     set_uxn_opcodes_phased_h_l353_c3_8c81_add <= VAR_set_uxn_opcodes_phased_h_l353_c3_8c81_add;
     -- Outputs

     -- t8_MUX[uxn_opcodes_phased_h_l343_c7_b0dd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond;
     t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output := t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l349_c7_789d] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond;
     result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue;
     result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output := result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l358_c7_d34c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l349_c7_789d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_cond;
     n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output := n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l355_c1_06d3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output;

     -- Submodule level 7
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c7_d34c_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l355_c1_06d3_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l349_c7_789d_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l346_c7_d915] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond;
     n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output := n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;

     -- put_stack[uxn_opcodes_phased_h_l356_c3_adfd] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l356_c3_adfd_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l356_c3_adfd_sp <= VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_sp;
     put_stack_uxn_opcodes_phased_h_l356_c3_adfd_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_stack_index;
     put_stack_uxn_opcodes_phased_h_l356_c3_adfd_offset <= VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_offset;
     put_stack_uxn_opcodes_phased_h_l356_c3_adfd_value <= VAR_put_stack_uxn_opcodes_phased_h_l356_c3_adfd_value;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l358_c1_f6de] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l346_c7_d915] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_cond;
     result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iftrue;
     result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output := result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l361_c7_6668] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l340_c2_b15f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond;
     t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output := t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;

     -- Submodule level 8
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c7_6668_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l358_c1_f6de_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l346_c7_d915_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;
     -- put_stack[uxn_opcodes_phased_h_l359_c3_2fb0] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_sp <= VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_sp;
     put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_stack_index;
     put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_offset <= VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_offset;
     put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_value <= VAR_put_stack_uxn_opcodes_phased_h_l359_c3_2fb0_value;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l361_c1_8ca3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l343_c7_b0dd] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond;
     result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue;
     result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output := result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l343_c7_b0dd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_cond;
     n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output := n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;

     -- Submodule level 9
     VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l361_c1_8ca3_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l343_c7_b0dd_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l340_c2_b15f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond;
     n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output := n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l340_c2_b15f] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_cond;
     result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iftrue;
     result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output := result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;

     -- put_stack[uxn_opcodes_phased_h_l362_c3_9e5b] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_sp <= VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_sp;
     put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_stack_index;
     put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_offset <= VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_offset;
     put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_value <= VAR_put_stack_uxn_opcodes_phased_h_l362_c3_9e5b_value;
     -- Outputs

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l340_c2_b15f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
