-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity ldz_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_f74745d5;
architecture arch of ldz_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1369_c6_1222]
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1369_c1_49f4]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal t8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1369_c2_31f8]
signal tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1370_c3_2262[uxn_opcodes_h_l1370_c3_2262]
signal printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1374_c11_1fb1]
signal BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal t8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1374_c7_74ae]
signal tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1377_c11_400b]
signal BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal t8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1377_c7_1e04]
signal tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1380_c30_3df1]
signal sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1383_c11_cb8c]
signal BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1383_c7_1142]
signal result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1383_c7_1142]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1383_c7_1142]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1383_c7_1142]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1383_c7_1142]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1383_c7_1142]
signal tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1386_c11_630a]
signal BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1386_c7_bdbe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1386_c7_bdbe]
signal result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1386_c7_bdbe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1386_c7_bdbe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1386_c7_bdbe]
signal tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1392_c11_da49]
signal BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1392_c7_b94d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1392_c7_b94d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a310( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222
BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_left,
BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_right,
BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output);

-- t8_MUX_uxn_opcodes_h_l1369_c2_31f8
t8_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8
result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8
result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8
tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond,
tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue,
tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse,
tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

-- printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262
printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262 : entity work.printf_uxn_opcodes_h_l1370_c3_2262_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1
BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_left,
BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_right,
BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output);

-- t8_MUX_uxn_opcodes_h_l1374_c7_74ae
t8_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae
result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae
result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae
result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae
result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae
result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae
result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae
tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond,
tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue,
tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse,
tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b
BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_left,
BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_right,
BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output);

-- t8_MUX_uxn_opcodes_h_l1377_c7_1e04
t8_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04
result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04
result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04
result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04
result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04
result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04
result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04
tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond,
tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue,
tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse,
tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1
sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_ins,
sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_x,
sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_y,
sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c
BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_left,
BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_right,
BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142
result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_cond,
result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142
result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142
result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142
result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1383_c7_1142
tmp8_MUX_uxn_opcodes_h_l1383_c7_1142 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_cond,
tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue,
tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse,
tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a
BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_left,
BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_right,
BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe
result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond,
result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe
result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe
result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe
tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond,
tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue,
tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse,
tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49
BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_left,
BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_right,
BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d
result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d
result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output,
 t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output,
 t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output,
 t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output,
 sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output,
 tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output,
 tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1371_c3_8a28 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_8c41 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1381_c22_02cc_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1389_c3_02ab : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_94d7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1369_l1383_l1374_DUPLICATE_1250_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_948a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1383_l1386_l1377_DUPLICATE_53d4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1397_l1365_DUPLICATE_daee_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1371_c3_8a28 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1371_c3_8a28;
     VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_8c41 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_8c41;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1389_c3_02ab := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1389_c3_02ab;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1383_c11_cb8c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_948a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_948a_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1381_c22_02cc] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1381_c22_02cc_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1377_c11_400b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1369_l1383_l1374_DUPLICATE_1250 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1369_l1383_l1374_DUPLICATE_1250_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1383_l1386_l1377_DUPLICATE_53d4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1383_l1386_l1377_DUPLICATE_53d4_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1374_c11_1fb1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1369_c6_1222] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_left;
     BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output := BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1392_c11_da49] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_left;
     BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output := BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1386_c11_630a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1380_c30_3df1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_ins;
     sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_x;
     sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output := sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output := result.u8_value;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_94d7 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_94d7_return_output := result.u16_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c6_1222_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1374_c11_1fb1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1377_c11_400b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1383_c11_cb8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1386_c11_630a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1392_c11_da49_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1381_c22_02cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_948a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_948a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_948a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_94d7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_94d7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1369_l1374_l1377_DUPLICATE_94d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1392_l1386_l1383_l1377_l1374_DUPLICATE_d7fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1369_l1383_l1374_DUPLICATE_1250_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1369_l1383_l1374_DUPLICATE_1250_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1369_l1383_l1374_DUPLICATE_1250_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1369_l1392_l1383_l1377_l1374_DUPLICATE_5d5c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1383_l1386_l1377_DUPLICATE_53d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1383_l1386_l1377_DUPLICATE_53d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1383_l1386_l1377_DUPLICATE_53d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1369_l1386_l1383_l1377_l1374_DUPLICATE_2f7c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1380_c30_3df1_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1386_c7_bdbe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output := result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;

     -- t8_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1386_c7_bdbe] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond;
     tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output := tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1386_c7_bdbe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1392_c7_b94d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1392_c7_b94d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1369_c1_49f4] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1383_c7_1142] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1369_c1_49f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1392_c7_b94d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1386_c7_bdbe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1383_c7_1142] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_cond;
     tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output := tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1383_c7_1142] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1386_c7_bdbe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;

     -- t8_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- printf_uxn_opcodes_h_l1370_c3_2262[uxn_opcodes_h_l1370_c3_2262] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1370_c3_2262_uxn_opcodes_h_l1370_c3_2262_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1383_c7_1142] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output := result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1386_c7_bdbe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1383_c7_1142] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- t8_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1383_c7_1142] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1383_c7_1142_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1377_c7_1e04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1377_c7_1e04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1374_c7_74ae] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1374_c7_74ae_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1369_c2_31f8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1397_l1365_DUPLICATE_daee LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1397_l1365_DUPLICATE_daee_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a310(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c2_31f8_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1397_l1365_DUPLICATE_daee_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1397_l1365_DUPLICATE_daee_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
