-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 64
entity sta2_0CLK_4674db74 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta2_0CLK_4674db74;
architecture arch of sta2_0CLK_4674db74 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_n16_high : unsigned(7 downto 0);
signal REG_COMB_n16_low : unsigned(7 downto 0);
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2339_c6_ccde]
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal t16_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(15 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2339_c2_2d30]
signal n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2352_c11_d501]
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal t16_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(15 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2352_c7_ce73]
signal n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2355_c11_63de]
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2355_c7_e098]
signal t16_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(15 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2355_c7_e098]
signal n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2355_c7_e098]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2355_c7_e098]
signal result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2355_c7_e098]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2355_c7_e098]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2355_c7_e098]
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2355_c7_e098]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2355_c7_e098]
signal n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2357_c3_8686]
signal CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2360_c11_6d04]
signal BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(15 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2360_c7_ea9c]
signal n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2361_c3_445a]
signal BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2364_c11_ef52]
signal BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(7 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2364_c7_8c33]
signal n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2366_c30_acc4]
signal sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2371_c11_f299]
signal BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2371_c7_b629]
signal result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2371_c7_b629]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2371_c7_b629]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2371_c7_b629]
signal result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(7 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2371_c7_b629]
signal n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l2374_c22_edc0]
signal BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output : unsigned(16 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_6145( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.is_stack_index_flipped := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;
      base.stack_address_sp_offset := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde
BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_left,
BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_right,
BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output);

-- t16_MUX_uxn_opcodes_h_l2339_c2_2d30
t16_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30
n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30
result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30
result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30
result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30
result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30
n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_cond,
n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue,
n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse,
n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_left,
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_right,
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output);

-- t16_MUX_uxn_opcodes_h_l2352_c7_ce73
t16_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73
n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73
result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73
result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73
n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_cond,
n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue,
n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse,
n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_left,
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_right,
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output);

-- t16_MUX_uxn_opcodes_h_l2355_c7_e098
t16_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
t16_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
t16_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2355_c7_e098
n16_high_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098
result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098
result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2355_c7_e098
n16_low_MUX_uxn_opcodes_h_l2355_c7_e098 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_cond,
n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue,
n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse,
n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2357_c3_8686
CONST_SL_8_uxn_opcodes_h_l2357_c3_8686 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_x,
CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_left,
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_right,
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output);

-- t16_MUX_uxn_opcodes_h_l2360_c7_ea9c
t16_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c
n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c
result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c
result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c
n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond,
n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue,
n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse,
n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a
BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_left,
BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_right,
BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52
BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_left,
BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_right,
BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33
n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33
result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33
result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33
result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33
result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33
result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33
n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_cond,
n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue,
n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse,
n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4
sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_ins,
sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_x,
sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_y,
sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299
BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_left,
BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_right,
BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629
result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond,
result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629
result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629
result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629
result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond,
result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2371_c7_b629
n16_low_MUX_uxn_opcodes_h_l2371_c7_b629 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_cond,
n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue,
n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse,
n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0
BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_left,
BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_right,
BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 n16_high,
 n16_low,
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output,
 t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output,
 t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output,
 t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output,
 CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output,
 t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output,
 n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output,
 sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output,
 n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2344_c3_5b78 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_0df3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2353_c3_9915 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2358_c3_7fc4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2362_c3_0c15 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_c7_ea9c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l2374_c3_9956 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2373_c3_3dbd : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output : unsigned(16 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2356_l2361_DUPLICATE_7b32_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l2379_l2334_DUPLICATE_d711_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_n16_high : unsigned(7 downto 0);
variable REG_VAR_n16_low : unsigned(7 downto 0);
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n16_high := n16_high;
  REG_VAR_n16_low := n16_low;
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_y := to_signed(-4, 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2344_c3_5b78 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2344_c3_5b78;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2358_c3_7fc4 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2358_c3_7fc4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2353_c3_9915 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2353_c3_9915;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_0df3 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_0df3;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2373_c3_3dbd := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2373_c3_3dbd;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2362_c3_0c15 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2362_c3_0c15;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_right := to_unsigned(5, 3);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_ins := VAR_ins;
     VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := n16_high;
     VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse := n16_low;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_left := VAR_phase;
     VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := VAR_previous_stack_read;
     VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_left := t16;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := t16;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2352_c11_d501] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_left;
     BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output := BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2339_c6_ccde] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_left;
     BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output := BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2366_c30_acc4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_ins;
     sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_x;
     sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output := sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l2374_c22_edc0] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_left;
     BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output := BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2356_l2361_DUPLICATE_7b32 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2356_l2361_DUPLICATE_7b32_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2364_c11_ef52] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_left;
     BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output := BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output := result.u16_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2355_c11_63de] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_left;
     BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output := BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2360_c11_6d04] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_left;
     BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output := BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_c7_ea9c_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2371_c11_f299] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_left;
     BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output := BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output;

     -- Submodule level 1
     VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c6_ccde_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_d501_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_63de_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_6d04_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2364_c11_ef52_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2371_c11_f299_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l2374_c3_9956 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l2374_c22_edc0_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2356_l2361_DUPLICATE_7b32_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2356_l2361_DUPLICATE_7b32_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2355_l2352_l2371_l2360_DUPLICATE_73ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_cda8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2371_l2364_l2360_l2355_DUPLICATE_883f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2364_l2355_l2352_l2360_DUPLICATE_05c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2352_l2339_l2371_l2360_l2355_DUPLICATE_1f37_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2339_c2_2d30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2366_c30_acc4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue := VAR_result_u16_value_uxn_opcodes_h_l2374_c3_9956;
     -- n16_low_MUX[uxn_opcodes_h_l2371_c7_b629] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_cond;
     n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output := n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2371_c7_b629] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output := result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2371_c7_b629] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2371_c7_b629] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2357_c3_8686] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output := CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2371_c7_b629] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output := result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2361_c3_445a] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_left;
     BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output := BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2361_c3_445a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2357_c3_8686_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2371_c7_b629_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- t16_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2364_c7_8c33] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- Submodule level 3
     VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2364_c7_8c33_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     -- n16_high_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2360_c7_ea9c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;

     -- t16_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     t16_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     t16_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- Submodule level 4
     VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_ea9c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2355_c7_e098] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output := result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;

     -- t16_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- Submodule level 5
     VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_e098_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2352_c7_ce73] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;

     -- t16_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- Submodule level 6
     REG_VAR_n16_high := VAR_n16_high_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_ce73_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2339_c2_2d30] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output := result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;

     -- Submodule level 7
     REG_VAR_n16_low := VAR_n16_low_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l2379_l2334_DUPLICATE_d711 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l2379_l2334_DUPLICATE_d711_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_6145(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2339_c2_2d30_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l2379_l2334_DUPLICATE_d711_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l2379_l2334_DUPLICATE_d711_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n16_high <= REG_VAR_n16_high;
REG_COMB_n16_low <= REG_VAR_n16_low;
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n16_high <= REG_COMB_n16_high;
     n16_low <= REG_COMB_n16_low;
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
