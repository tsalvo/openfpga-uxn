-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 7
entity opc_dup_0CLK_908f9b38 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_dup_0CLK_908f9b38;
architecture arch of opc_dup_0CLK_908f9b38 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- t_register[uxn_opcodes_h_l214_c7_69e7]
signal t_register_uxn_opcodes_h_l214_c7_69e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_h_l214_c7_69e7_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_h_l214_c7_69e7_return_output : unsigned(7 downto 0);

-- set[uxn_opcodes_h_l215_c9_43ee]
signal set_uxn_opcodes_h_l215_c9_43ee_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_h_l215_c9_43ee_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_h_l215_c9_43ee_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_h_l215_c9_43ee_k : unsigned(7 downto 0);
signal set_uxn_opcodes_h_l215_c9_43ee_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_h_l215_c9_43ee_add : signed(7 downto 0);
signal set_uxn_opcodes_h_l215_c9_43ee_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l216_c6_4cff]
signal BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l217_c1_2eaa]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_h_l216_c2_4676]
signal result_MUX_uxn_opcodes_h_l216_c2_4676_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l216_c2_4676_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l216_c2_4676_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l216_c2_4676_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_h_l218_c3_0f0c]
signal put_stack_uxn_opcodes_h_l218_c3_0f0c_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_h_l218_c3_0f0c_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_h_l218_c3_0f0c_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_h_l218_c3_0f0c_value : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_h_l219_c3_777c]
signal put_stack_uxn_opcodes_h_l219_c3_777c_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_h_l219_c3_777c_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_h_l219_c3_777c_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_h_l219_c3_777c_value : unsigned(7 downto 0);


begin

-- SUBMODULE INSTANCES 
-- t_register_uxn_opcodes_h_l214_c7_69e7
t_register_uxn_opcodes_h_l214_c7_69e7 : entity work.t_register_0CLK_0e5af5c0 port map (
clk,
t_register_uxn_opcodes_h_l214_c7_69e7_CLOCK_ENABLE,
t_register_uxn_opcodes_h_l214_c7_69e7_stack_index,
t_register_uxn_opcodes_h_l214_c7_69e7_return_output);

-- set_uxn_opcodes_h_l215_c9_43ee
set_uxn_opcodes_h_l215_c9_43ee : entity work.set_0CLK_e105ce74 port map (
clk,
set_uxn_opcodes_h_l215_c9_43ee_CLOCK_ENABLE,
set_uxn_opcodes_h_l215_c9_43ee_stack_index,
set_uxn_opcodes_h_l215_c9_43ee_ins,
set_uxn_opcodes_h_l215_c9_43ee_k,
set_uxn_opcodes_h_l215_c9_43ee_mul,
set_uxn_opcodes_h_l215_c9_43ee_add,
set_uxn_opcodes_h_l215_c9_43ee_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff
BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_left,
BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_right,
BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output);

-- result_MUX_uxn_opcodes_h_l216_c2_4676
result_MUX_uxn_opcodes_h_l216_c2_4676 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_h_l216_c2_4676_cond,
result_MUX_uxn_opcodes_h_l216_c2_4676_iftrue,
result_MUX_uxn_opcodes_h_l216_c2_4676_iffalse,
result_MUX_uxn_opcodes_h_l216_c2_4676_return_output);

-- put_stack_uxn_opcodes_h_l218_c3_0f0c
put_stack_uxn_opcodes_h_l218_c3_0f0c : entity work.put_stack_0CLK_e3ba3c7d port map (
clk,
put_stack_uxn_opcodes_h_l218_c3_0f0c_CLOCK_ENABLE,
put_stack_uxn_opcodes_h_l218_c3_0f0c_stack_index,
put_stack_uxn_opcodes_h_l218_c3_0f0c_offset,
put_stack_uxn_opcodes_h_l218_c3_0f0c_value);

-- put_stack_uxn_opcodes_h_l219_c3_777c
put_stack_uxn_opcodes_h_l219_c3_777c : entity work.put_stack_0CLK_e3ba3c7d port map (
clk,
put_stack_uxn_opcodes_h_l219_c3_777c_CLOCK_ENABLE,
put_stack_uxn_opcodes_h_l219_c3_777c_stack_index,
put_stack_uxn_opcodes_h_l219_c3_777c_offset,
put_stack_uxn_opcodes_h_l219_c3_777c_value);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 stack_index,
 ins,
 k,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 t_register_uxn_opcodes_h_l214_c7_69e7_return_output,
 set_uxn_opcodes_h_l215_c9_43ee_return_output,
 BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output,
 result_MUX_uxn_opcodes_h_l216_c2_4676_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_h_l214_c7_69e7_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_h_l214_c7_69e7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_h_l214_c7_69e7_return_output : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_h_l215_c9_43ee_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l219_c3_777c_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l219_c3_777c_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l219_c3_777c_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_h_l219_c3_777c_CLOCK_ENABLE : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_put_stack_uxn_opcodes_h_l219_c3_777c_offset := resize(to_unsigned(1, 1), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iftrue := to_unsigned(0, 1);
     VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_offset := resize(to_unsigned(0, 1), 8);
     VAR_set_uxn_opcodes_h_l215_c9_43ee_mul := resize(to_unsigned(1, 1), 8);
     VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_iftrue := to_unsigned(1, 1);
     VAR_set_uxn_opcodes_h_l215_c9_43ee_add := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iffalse := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_h_l215_c9_43ee_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_t_register_uxn_opcodes_h_l214_c7_69e7_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_h_l215_c9_43ee_ins := VAR_ins;
     VAR_set_uxn_opcodes_h_l215_c9_43ee_k := VAR_k;
     VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_h_l219_c3_777c_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_h_l215_c9_43ee_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_h_l214_c7_69e7_stack_index := VAR_stack_index;
     -- set[uxn_opcodes_h_l215_c9_43ee] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_h_l215_c9_43ee_CLOCK_ENABLE <= VAR_set_uxn_opcodes_h_l215_c9_43ee_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_h_l215_c9_43ee_stack_index <= VAR_set_uxn_opcodes_h_l215_c9_43ee_stack_index;
     set_uxn_opcodes_h_l215_c9_43ee_ins <= VAR_set_uxn_opcodes_h_l215_c9_43ee_ins;
     set_uxn_opcodes_h_l215_c9_43ee_k <= VAR_set_uxn_opcodes_h_l215_c9_43ee_k;
     set_uxn_opcodes_h_l215_c9_43ee_mul <= VAR_set_uxn_opcodes_h_l215_c9_43ee_mul;
     set_uxn_opcodes_h_l215_c9_43ee_add <= VAR_set_uxn_opcodes_h_l215_c9_43ee_add;
     -- Outputs
     VAR_set_uxn_opcodes_h_l215_c9_43ee_return_output := set_uxn_opcodes_h_l215_c9_43ee_return_output;

     -- t_register[uxn_opcodes_h_l214_c7_69e7] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_h_l214_c7_69e7_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_h_l214_c7_69e7_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_h_l214_c7_69e7_stack_index <= VAR_t_register_uxn_opcodes_h_l214_c7_69e7_stack_index;
     -- Outputs
     VAR_t_register_uxn_opcodes_h_l214_c7_69e7_return_output := t_register_uxn_opcodes_h_l214_c7_69e7_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_left := VAR_set_uxn_opcodes_h_l215_c9_43ee_return_output;
     REG_VAR_tmp8 := VAR_set_uxn_opcodes_h_l215_c9_43ee_return_output;
     VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_value := VAR_t_register_uxn_opcodes_h_l214_c7_69e7_return_output;
     VAR_put_stack_uxn_opcodes_h_l219_c3_777c_value := VAR_t_register_uxn_opcodes_h_l214_c7_69e7_return_output;
     REG_VAR_t8 := VAR_t_register_uxn_opcodes_h_l214_c7_69e7_return_output;
     -- BIN_OP_GT[uxn_opcodes_h_l216_c6_4cff] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_left;
     BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output := BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output;
     VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l216_c6_4cff_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l217_c1_2eaa] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output;

     -- result_MUX[uxn_opcodes_h_l216_c2_4676] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_h_l216_c2_4676_cond <= VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_cond;
     result_MUX_uxn_opcodes_h_l216_c2_4676_iftrue <= VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_iftrue;
     result_MUX_uxn_opcodes_h_l216_c2_4676_iffalse <= VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_return_output := result_MUX_uxn_opcodes_h_l216_c2_4676_return_output;

     -- Submodule level 3
     VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output;
     VAR_put_stack_uxn_opcodes_h_l219_c3_777c_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l217_c1_2eaa_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_h_l216_c2_4676_return_output;
     -- put_stack[uxn_opcodes_h_l219_c3_777c] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_h_l219_c3_777c_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_h_l219_c3_777c_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_h_l219_c3_777c_stack_index <= VAR_put_stack_uxn_opcodes_h_l219_c3_777c_stack_index;
     put_stack_uxn_opcodes_h_l219_c3_777c_offset <= VAR_put_stack_uxn_opcodes_h_l219_c3_777c_offset;
     put_stack_uxn_opcodes_h_l219_c3_777c_value <= VAR_put_stack_uxn_opcodes_h_l219_c3_777c_value;
     -- Outputs

     -- put_stack[uxn_opcodes_h_l218_c3_0f0c] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_h_l218_c3_0f0c_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_h_l218_c3_0f0c_stack_index <= VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_stack_index;
     put_stack_uxn_opcodes_h_l218_c3_0f0c_offset <= VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_offset;
     put_stack_uxn_opcodes_h_l218_c3_0f0c_value <= VAR_put_stack_uxn_opcodes_h_l218_c3_0f0c_value;
     -- Outputs

     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
