-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity dup2_0CLK_3554410e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup2_0CLK_3554410e;
architecture arch of dup2_0CLK_3554410e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2751_c6_713a]
signal BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2751_c2_4c41]
signal t16_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2751_c2_4c41]
signal result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2751_c2_4c41]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2751_c2_4c41]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2751_c2_4c41]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2751_c2_4c41]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2758_c11_d5ad]
signal BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2758_c7_8280]
signal t16_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2758_c7_8280]
signal result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2758_c7_8280]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2758_c7_8280]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2758_c7_8280]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2758_c7_8280]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2761_c11_1414]
signal BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2761_c7_512e]
signal t16_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2761_c7_512e]
signal result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2761_c7_512e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2761_c7_512e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2761_c7_512e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2761_c7_512e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2763_c3_3a34]
signal CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2765_c30_b205]
signal sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2767_c11_c195]
signal BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2767_c7_9397]
signal t16_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2767_c7_9397]
signal result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2767_c7_9397]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2767_c7_9397]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2767_c7_9397]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2767_c7_9397]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2768_c3_eba6]
signal BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2774_c11_73f5]
signal BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2774_c7_7987]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2774_c7_7987]
signal result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2774_c7_7987]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2774_c7_7987]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2778_c11_8df6]
signal BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2778_c7_c346]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2778_c7_c346]
signal result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2778_c7_c346]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2778_c7_c346]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2782_c11_d560]
signal BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2782_c7_2a1e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2782_c7_2a1e]
signal result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2782_c7_2a1e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2782_c7_2a1e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2786_c11_b60a]
signal BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2786_c7_7496]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2786_c7_7496]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output : unsigned(0 downto 0);

-- CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6
signal CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_x : unsigned(15 downto 0);
signal CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output : unsigned(15 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a
BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_left,
BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_right,
BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output);

-- t16_MUX_uxn_opcodes_h_l2751_c2_4c41
t16_MUX_uxn_opcodes_h_l2751_c2_4c41 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2751_c2_4c41_cond,
t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue,
t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse,
t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41
result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_cond,
result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41
result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41
result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41
result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad
BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_left,
BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_right,
BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output);

-- t16_MUX_uxn_opcodes_h_l2758_c7_8280
t16_MUX_uxn_opcodes_h_l2758_c7_8280 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2758_c7_8280_cond,
t16_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue,
t16_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse,
t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280
result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_cond,
result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280
result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280
result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280
result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414
BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_left,
BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_right,
BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output);

-- t16_MUX_uxn_opcodes_h_l2761_c7_512e
t16_MUX_uxn_opcodes_h_l2761_c7_512e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2761_c7_512e_cond,
t16_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue,
t16_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse,
t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e
result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e
result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e
result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34
CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_x,
CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2765_c30_b205
sp_relative_shift_uxn_opcodes_h_l2765_c30_b205 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_ins,
sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_x,
sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_y,
sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195
BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_left,
BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_right,
BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output);

-- t16_MUX_uxn_opcodes_h_l2767_c7_9397
t16_MUX_uxn_opcodes_h_l2767_c7_9397 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2767_c7_9397_cond,
t16_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue,
t16_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse,
t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397
result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_cond,
result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397
result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397
result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397
result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6
BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_left,
BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_right,
BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5
BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_left,
BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_right,
BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987
result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987
result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_cond,
result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987
result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6
BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_left,
BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_right,
BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346
result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346
result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_cond,
result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346
result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560
BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_left,
BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_right,
BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e
result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e
result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e
result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_left,
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_right,
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output);

-- CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6
CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_x,
CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output,
 t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output,
 t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output,
 t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output,
 CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output,
 sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output,
 t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output,
 CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2755_c3_962a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2759_c3_e111 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_x : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2771_c3_20f6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2769_c3_dc2f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2772_c21_4817_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2775_c3_5c0b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2779_c3_d433 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2780_c21_9328_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2783_c3_deed : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2751_l2767_l2758_DUPLICATE_770b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2762_l2768_DUPLICATE_08f9_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2761_l2782_DUPLICATE_8c98_return_output : unsigned(3 downto 0);
 variable VAR_CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_x : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uint16_t_uxn_opcodes_h_l2784_l2776_DUPLICATE_a9bb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2791_l2747_DUPLICATE_251e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_right := to_unsigned(6, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2759_c3_e111 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2759_c3_e111;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2771_c3_20f6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2771_c3_20f6;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2775_c3_5c0b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2775_c3_5c0b;
     VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2783_c3_deed := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2783_c3_deed;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2755_c3_962a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2755_c3_962a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2779_c3_d433 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2779_c3_d433;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_right := to_unsigned(4, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2769_c3_dc2f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2769_c3_dc2f;
     VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_left := t16;
     VAR_CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_x := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2778_c11_8df6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2762_l2768_DUPLICATE_08f9 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2762_l2768_DUPLICATE_08f9_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2761_l2782_DUPLICATE_8c98 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2761_l2782_DUPLICATE_8c98_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2761_c11_1414] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_left;
     BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output := BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2751_l2767_l2758_DUPLICATE_770b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2751_l2767_l2758_DUPLICATE_770b_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2758_c11_d5ad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_left;
     BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output := BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2786_c11_b60a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output;

     -- CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6 LATENCY=0
     -- Inputs
     CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_x <= VAR_CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_x;
     -- Outputs
     VAR_CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output := CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2751_c6_713a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2765_c30_b205] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_ins;
     sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_x;
     sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output := sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2767_c11_c195] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_left;
     BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output := BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2780_c21_9328] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2780_c21_9328_return_output := CAST_TO_uint8_t_uint16_t(
     t16);

     -- BIN_OP_EQ[uxn_opcodes_h_l2782_c11_d560] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_left;
     BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output := BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2774_c11_73f5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2751_c6_713a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2758_c11_d5ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2761_c11_1414_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2767_c11_c195_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2774_c11_73f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2778_c11_8df6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2782_c11_d560_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_b60a_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2762_l2768_DUPLICATE_08f9_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2762_l2768_DUPLICATE_08f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2780_c21_9328_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2751_l2767_l2758_DUPLICATE_770b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2751_l2767_l2758_DUPLICATE_770b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2751_l2767_l2758_DUPLICATE_770b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2774_l2767_l2761_l2758_l2786_l2782_l2778_DUPLICATE_f078_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2774_l2761_l2758_l2786_l2751_l2782_l2778_DUPLICATE_bbec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2761_l2782_DUPLICATE_8c98_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2761_l2782_DUPLICATE_8c98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2761_l2751_l2782_l2758_DUPLICATE_35bf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2765_c30_b205_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2767_c7_9397] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2768_c3_eba6] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_left;
     BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output := BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2763_c3_3a34] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output := CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2786_c7_7496] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2786_c7_7496] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output;

     -- CAST_TO_uint8_t_uint16_t_uxn_opcodes_h_l2784_l2776_DUPLICATE_a9bb LATENCY=0
     VAR_CAST_TO_uint8_t_uint16_t_uxn_opcodes_h_l2784_l2776_DUPLICATE_a9bb_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uint16_t_uxn_opcodes_h_l2776_l2784_DUPLICATE_dcb6_return_output);

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2782_c7_2a1e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue := VAR_CAST_TO_uint8_t_uint16_t_uxn_opcodes_h_l2784_l2776_DUPLICATE_a9bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue := VAR_CAST_TO_uint8_t_uint16_t_uxn_opcodes_h_l2784_l2776_DUPLICATE_a9bb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2763_c3_3a34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_7496_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_7496_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;
     -- CAST_TO_uint8_t[uxn_opcodes_h_l2772_c21_4817] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2772_c21_4817_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l2768_c3_eba6_return_output);

     -- result_u8_value_MUX[uxn_opcodes_h_l2782_c7_2a1e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2761_c7_512e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;

     -- t16_MUX[uxn_opcodes_h_l2767_c7_9397] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2767_c7_9397_cond <= VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_cond;
     t16_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue;
     t16_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output := t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2782_c7_2a1e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2782_c7_2a1e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2778_c7_c346] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2772_c21_4817_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2782_c7_2a1e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;
     -- t16_MUX[uxn_opcodes_h_l2761_c7_512e] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2761_c7_512e_cond <= VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_cond;
     t16_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue;
     t16_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output := t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2758_c7_8280] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2778_c7_c346] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2774_c7_7987] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2778_c7_c346] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2778_c7_c346] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output := result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2778_c7_c346_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2751_c2_4c41] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;

     -- t16_MUX[uxn_opcodes_h_l2758_c7_8280] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2758_c7_8280_cond <= VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_cond;
     t16_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue;
     t16_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output := t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2767_c7_9397] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2774_c7_7987] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output := result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2774_c7_7987] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2774_c7_7987] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2774_c7_7987_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2761_c7_512e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;

     -- t16_MUX[uxn_opcodes_h_l2751_c2_4c41] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2751_c2_4c41_cond <= VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_cond;
     t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue;
     t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output := t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2767_c7_9397] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2767_c7_9397] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2767_c7_9397] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output := result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2767_c7_9397_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2758_c7_8280] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2761_c7_512e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2761_c7_512e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2761_c7_512e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2761_c7_512e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2758_c7_8280] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2751_c2_4c41] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2758_c7_8280] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output := result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2758_c7_8280] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;

     -- Submodule level 8
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2758_c7_8280_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2751_c2_4c41] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2751_c2_4c41] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output := result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2751_c2_4c41] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2791_l2747_DUPLICATE_251e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2791_l2747_DUPLICATE_251e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2751_c2_4c41_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2791_l2747_DUPLICATE_251e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2791_l2747_DUPLICATE_251e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
