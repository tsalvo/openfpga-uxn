-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity deo_0CLK_da9cb8d4 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 previous_device_ram_read : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end deo_0CLK_da9cb8d4;
architecture arch of deo_0CLK_da9cb8d4 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal device_out_result : device_out_result_t := device_out_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;
signal REG_COMB_device_out_result : device_out_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l483_c6_2ab8]
signal BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l491_c7_9d67]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_is_device_ram_16bit_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(15 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(23 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(23 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(23 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l483_c2_a182]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l483_c2_a182]
signal t8_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l483_c2_a182]
signal n8_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l483_c2_a182]
signal device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output : device_out_result_t;

-- BIN_OP_EQ[uxn_opcodes_h_l491_c11_d670]
signal BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l496_c1_a162]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output : unsigned(0 downto 0);

-- result_is_device_ram_16bit_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : signed(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(23 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(23 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(23 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l491_c7_9d67]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l491_c7_9d67]
signal t8_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l491_c7_9d67]
signal n8_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l491_c7_9d67]
signal device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : device_out_result_t;

-- sp_relative_shift[uxn_opcodes_h_l494_c30_51e6]
signal sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l497_c9_51dc]
signal BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l497_c9_b6c1]
signal MUX_uxn_opcodes_h_l497_c9_b6c1_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l497_c9_b6c1_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l497_c9_b6c1_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l497_c9_b6c1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l498_c9_4031]
signal BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l498_c33_79d3]
signal CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output : unsigned(15 downto 0);

-- MUX[uxn_opcodes_h_l498_c9_a42d]
signal MUX_uxn_opcodes_h_l498_c9_a42d_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l498_c9_a42d_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l498_c9_a42d_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l498_c9_a42d_return_output : unsigned(7 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l500_c42_fbcc]
signal BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output : unsigned(7 downto 0);

-- device_out[uxn_opcodes_h_l500_c23_29d4]
signal device_out_uxn_opcodes_h_l500_c23_29d4_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_out_uxn_opcodes_h_l500_c23_29d4_device_address : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l500_c23_29d4_value : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l500_c23_29d4_phase : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l500_c23_29d4_previous_device_ram_read : unsigned(15 downto 0);
signal device_out_uxn_opcodes_h_l500_c23_29d4_previous_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l500_c23_29d4_return_output : device_out_result_t;

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_aff6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_device_ram_16bit := ref_toks_1;
      base.device_ram_address := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_device_ram_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;
      base.vram_write_layer := ref_toks_10;
      base.vram_address := ref_toks_11;
      base.is_sp_shift := ref_toks_12;
      base.is_stack_operation_16bit := ref_toks_13;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8
BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_left,
BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_right,
BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182
result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182
result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182
result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182
result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182
result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182
result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182
result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182
result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182
result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint24_t_uint24_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182
result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- t8_MUX_uxn_opcodes_h_l483_c2_a182
t8_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l483_c2_a182_cond,
t8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
t8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- n8_MUX_uxn_opcodes_h_l483_c2_a182
n8_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l483_c2_a182_cond,
n8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
n8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l483_c2_a182
device_out_result_MUX_uxn_opcodes_h_l483_c2_a182 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_cond,
device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iftrue,
device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iffalse,
device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670
BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_left,
BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_right,
BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output);

-- result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67
result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67
result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67
result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67
result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67
result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67
result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67
result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67
result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67
result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint24_t_uint24_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67
result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- t8_MUX_uxn_opcodes_h_l491_c7_9d67
t8_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
t8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
t8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- n8_MUX_uxn_opcodes_h_l491_c7_9d67
n8_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
n8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
n8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67
device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_cond,
device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue,
device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse,
device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output);

-- sp_relative_shift_uxn_opcodes_h_l494_c30_51e6
sp_relative_shift_uxn_opcodes_h_l494_c30_51e6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_ins,
sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_x,
sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_y,
sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc
BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_left,
BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_right,
BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output);

-- MUX_uxn_opcodes_h_l497_c9_b6c1
MUX_uxn_opcodes_h_l497_c9_b6c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l497_c9_b6c1_cond,
MUX_uxn_opcodes_h_l497_c9_b6c1_iftrue,
MUX_uxn_opcodes_h_l497_c9_b6c1_iffalse,
MUX_uxn_opcodes_h_l497_c9_b6c1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031
BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_left,
BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_right,
BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output);

-- CONST_SR_8_uxn_opcodes_h_l498_c33_79d3
CONST_SR_8_uxn_opcodes_h_l498_c33_79d3 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_x,
CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output);

-- MUX_uxn_opcodes_h_l498_c9_a42d
MUX_uxn_opcodes_h_l498_c9_a42d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l498_c9_a42d_cond,
MUX_uxn_opcodes_h_l498_c9_a42d_iftrue,
MUX_uxn_opcodes_h_l498_c9_a42d_iffalse,
MUX_uxn_opcodes_h_l498_c9_a42d_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc
BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_left,
BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_right,
BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output);

-- device_out_uxn_opcodes_h_l500_c23_29d4
device_out_uxn_opcodes_h_l500_c23_29d4 : entity work.device_out_0CLK_8af766d2 port map (
clk,
device_out_uxn_opcodes_h_l500_c23_29d4_CLOCK_ENABLE,
device_out_uxn_opcodes_h_l500_c23_29d4_device_address,
device_out_uxn_opcodes_h_l500_c23_29d4_value,
device_out_uxn_opcodes_h_l500_c23_29d4_phase,
device_out_uxn_opcodes_h_l500_c23_29d4_previous_device_ram_read,
device_out_uxn_opcodes_h_l500_c23_29d4_previous_ram_read,
device_out_uxn_opcodes_h_l500_c23_29d4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 previous_ram_read,
 -- Registers
 t8,
 n8,
 result,
 device_out_result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output,
 result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output,
 sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output,
 MUX_uxn_opcodes_h_l497_c9_b6c1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output,
 CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output,
 MUX_uxn_opcodes_h_l498_c9_a42d_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output,
 device_out_uxn_opcodes_h_l500_c23_29d4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_previous_device_ram_read : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l488_c3_991a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(23 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(23 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(23 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(23 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(23 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(23 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l491_c7_9d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_iffalse : unsigned(7 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l497_c23_d5b6_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l498_c9_a42d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l498_c9_a42d_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l498_c9_a42d_iffalse : unsigned(7 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l498_c23_f7cb_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l498_c9_a42d_return_output : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_device_address : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_value : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_phase : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_previous_device_ram_read : unsigned(15 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output : device_out_result_t;
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l501_c32_0f31_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l502_c32_5e39_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l503_c31_ec09_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l504_c21_6206_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_value_d41d_uxn_opcodes_h_l505_c22_c1a2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l506_c26_98c5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l507_c29_b499_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint24_t_device_out_result_t_vram_address_d41d_uxn_opcodes_h_l508_c25_16e4_return_output : unsigned(23 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l509_c24_9f96_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_ef07_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9170_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_3fb3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_6876_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_7c8b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_c48f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9f26_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_8627_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint24_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_04da_return_output : unsigned(23 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_aff6_uxn_opcodes_h_l512_l478_DUPLICATE_f8de_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
variable REG_VAR_device_out_result : device_out_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
  REG_VAR_device_out_result := device_out_result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l488_c3_991a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l488_c3_991a;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_right := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := device_out_result;
     VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_ins := VAR_ins;
     VAR_MUX_uxn_opcodes_h_l498_c9_a42d_iffalse := n8;
     VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_left := VAR_phase;
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_previous_ram_read := VAR_previous_ram_read;
     VAR_CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_x := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l497_c9_51dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_left;
     BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output := BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_6876 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_6876_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l494_c30_51e6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_ins;
     sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_x;
     sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output := sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_c48f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_c48f_return_output := result.u8_value;

     -- result_is_opc_done_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     VAR_result_is_opc_done_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l491_c7_9d67_return_output := result.is_opc_done;

     -- BIN_OP_MINUS[uxn_opcodes_h_l500_c42_fbcc] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_left;
     BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output := BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9170 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9170_return_output := result.device_ram_address;

     -- BIN_OP_EQ[uxn_opcodes_h_l483_c6_2ab8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_left;
     BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output := BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;

     -- CONST_REF_RD_uint24_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_04da LATENCY=0
     VAR_CONST_REF_RD_uint24_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_04da_return_output := result.vram_address;

     -- BIN_OP_EQ[uxn_opcodes_h_l491_c11_d670] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_left;
     BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output := BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_ef07 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_ef07_return_output := result.is_device_ram_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_8627 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_8627_return_output := result.vram_write_layer;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9f26 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9f26_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_7c8b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_7c8b_return_output := result.is_device_ram_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l483_c2_a182_return_output := result.stack_address_sp_offset;

     -- result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l491_c7_9d67_return_output := result.is_stack_operation_16bit;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l497_c23_d5b6] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l497_c23_d5b6_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l498_c9_4031] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_left;
     BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output := BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output;

     -- result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     VAR_result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l483_c2_a182_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_3fb3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_3fb3_return_output := result.is_vram_write;

     -- CONST_SR_8[uxn_opcodes_h_l498_c33_79d3] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_x <= VAR_CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output := CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l483_c6_2ab8_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l491_c11_d670_return_output;
     VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l497_c9_51dc_return_output;
     VAR_MUX_uxn_opcodes_h_l498_c9_a42d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l498_c9_4031_return_output;
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l500_c42_fbcc_return_output;
     VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l497_c23_d5b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9f26_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9f26_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_6876_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_6876_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_ef07_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_ef07_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_7c8b_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_7c8b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_3fb3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_3fb3_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_8627_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_8627_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint24_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_04da_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint24_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_04da_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9170_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_9170_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_c48f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l483_l491_DUPLICATE_c48f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_result_is_opc_done_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue := VAR_result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l483_c2_a182_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l483_c2_a182_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l494_c30_51e6_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l498_c23_f7cb] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l498_c23_f7cb_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l498_c33_79d3_return_output);

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- MUX[uxn_opcodes_h_l497_c9_b6c1] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l497_c9_b6c1_cond <= VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_cond;
     MUX_uxn_opcodes_h_l497_c9_b6c1_iftrue <= VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_iftrue;
     MUX_uxn_opcodes_h_l497_c9_b6c1_iffalse <= VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_return_output := MUX_uxn_opcodes_h_l497_c9_b6c1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l498_c9_a42d_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l498_c23_f7cb_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_device_address := VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_MUX_uxn_opcodes_h_l497_c9_b6c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     -- t8_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     t8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     t8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- MUX[uxn_opcodes_h_l498_c9_a42d] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l498_c9_a42d_cond <= VAR_MUX_uxn_opcodes_h_l498_c9_a42d_cond;
     MUX_uxn_opcodes_h_l498_c9_a42d_iftrue <= VAR_MUX_uxn_opcodes_h_l498_c9_a42d_iftrue;
     MUX_uxn_opcodes_h_l498_c9_a42d_iffalse <= VAR_MUX_uxn_opcodes_h_l498_c9_a42d_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l498_c9_a42d_return_output := MUX_uxn_opcodes_h_l498_c9_a42d_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l496_c1_a162] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- Submodule level 3
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l496_c1_a162_return_output;
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_value := VAR_MUX_uxn_opcodes_h_l498_c9_a42d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_MUX_uxn_opcodes_h_l498_c9_a42d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_t8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     -- device_out[uxn_opcodes_h_l500_c23_29d4] LATENCY=0
     -- Clock enable
     device_out_uxn_opcodes_h_l500_c23_29d4_CLOCK_ENABLE <= VAR_device_out_uxn_opcodes_h_l500_c23_29d4_CLOCK_ENABLE;
     -- Inputs
     device_out_uxn_opcodes_h_l500_c23_29d4_device_address <= VAR_device_out_uxn_opcodes_h_l500_c23_29d4_device_address;
     device_out_uxn_opcodes_h_l500_c23_29d4_value <= VAR_device_out_uxn_opcodes_h_l500_c23_29d4_value;
     device_out_uxn_opcodes_h_l500_c23_29d4_phase <= VAR_device_out_uxn_opcodes_h_l500_c23_29d4_phase;
     device_out_uxn_opcodes_h_l500_c23_29d4_previous_device_ram_read <= VAR_device_out_uxn_opcodes_h_l500_c23_29d4_previous_device_ram_read;
     device_out_uxn_opcodes_h_l500_c23_29d4_previous_ram_read <= VAR_device_out_uxn_opcodes_h_l500_c23_29d4_previous_ram_read;
     -- Outputs
     VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output := device_out_uxn_opcodes_h_l500_c23_29d4_return_output;

     -- t8_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     t8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     t8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output := t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- n8_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     n8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     n8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- Submodule level 4
     VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_n8_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l483_c2_a182_return_output;
     -- n8_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     n8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     n8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output := n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d[uxn_opcodes_h_l507_c29_b499] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l507_c29_b499_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.vram_write_layer;

     -- device_out_result_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d[uxn_opcodes_h_l503_c31_ec09] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l503_c31_ec09_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.device_ram_address;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l501_c32_0f31] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l501_c32_0f31_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.is_device_ram_write;

     -- CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d[uxn_opcodes_h_l504_c21_6206] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l504_c21_6206_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.u8_value;

     -- CONST_REF_RD_uint24_t_device_out_result_t_vram_address_d41d[uxn_opcodes_h_l508_c25_16e4] LATENCY=0
     VAR_CONST_REF_RD_uint24_t_device_out_result_t_vram_address_d41d_uxn_opcodes_h_l508_c25_16e4_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.vram_address;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d[uxn_opcodes_h_l506_c26_98c5] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l506_c26_98c5_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.is_vram_write;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d[uxn_opcodes_h_l509_c24_9f96] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l509_c24_9f96_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.is_deo_done;

     -- CONST_REF_RD_uint16_t_device_out_result_t_u16_value_d41d[uxn_opcodes_h_l505_c22_c1a2] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_value_d41d_uxn_opcodes_h_l505_c22_c1a2_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.u16_value;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_16bit_d41d[uxn_opcodes_h_l502_c32_5e39] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l502_c32_5e39_return_output := VAR_device_out_uxn_opcodes_h_l500_c23_29d4_return_output.is_device_ram_16bit;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_value_d41d_uxn_opcodes_h_l505_c22_c1a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l509_c24_9f96_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l502_c32_5e39_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l501_c32_0f31_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l506_c26_98c5_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l507_c29_b499_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint24_t_device_out_result_t_vram_address_d41d_uxn_opcodes_h_l508_c25_16e4_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l503_c31_ec09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l504_c21_6206_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l483_c2_a182_return_output;
     -- result_vram_address_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_is_device_ram_16bit_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output := device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l491_c7_9d67] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;

     -- Submodule level 6
     REG_VAR_device_out_result := VAR_device_out_result_MUX_uxn_opcodes_h_l483_c2_a182_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_vram_address_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l491_c7_9d67_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_is_device_ram_16bit_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_vram_address_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l483_c2_a182] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_aff6_uxn_opcodes_h_l512_l478_DUPLICATE_f8de LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_aff6_uxn_opcodes_h_l512_l478_DUPLICATE_f8de_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_aff6(
     result,
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_vram_address_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l483_c2_a182_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l483_c2_a182_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_aff6_uxn_opcodes_h_l512_l478_DUPLICATE_f8de_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_aff6_uxn_opcodes_h_l512_l478_DUPLICATE_f8de_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
REG_COMB_device_out_result <= REG_VAR_device_out_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
     device_out_result <= REG_COMB_device_out_result;
 end if;
 end if;
end process;

end arch;
