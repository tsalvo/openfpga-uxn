-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_8;
 var_dim_0 : in unsigned(2 downto 0);
 return_output : out uint8_t_array_8_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_060a( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return uint8_t_array_8_t is
 
  variable base : uint8_t_array_8_t; 
  variable return_output : uint8_t_array_8_t;
begin
      base.data(1) := ref_toks_0;
      base.data(7) := ref_toks_1;
      base.data(4) := ref_toks_2;
      base.data(0) := ref_toks_3;
      base.data(3) := ref_toks_4;
      base.data(6) := ref_toks_5;
      base.data(2) := ref_toks_6;
      base.data(5) := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38 : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_8;
 variable VAR_var_dim_0 : unsigned(2 downto 0);
 variable VAR_return_output : uint8_t_array_8_t;
 variable VAR_base : uint8_t_8;
 variable VAR_rv : uint8_t_array_8_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_43e5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_4dbd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_4430_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_e8f9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_6ce3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_08fd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_0215_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_a975_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_060a_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_3347_return_output : uint8_t_array_8_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_a975] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_a975_return_output := VAR_ref_toks_0(5);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_6ce3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_6ce3_return_output := VAR_ref_toks_0(3);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_0215] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_0215_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_8_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_08fd] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_08fd_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_8_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_4430] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_4430_return_output := VAR_ref_toks_0(4);

     -- CONST_REF_RD_uint8_t_uint8_t_8_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_43e5] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_43e5_return_output := VAR_ref_toks_0(1);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_e8f9] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_e8f9_return_output := VAR_ref_toks_0(0);

     -- CONST_REF_RD_uint8_t_uint8_t_8_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_4dbd] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_4dbd_return_output := VAR_ref_toks_0(7);

     -- Submodule level 1
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_2e38_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_d03d_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_1d33_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_e9ba_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_e9da_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_9cac_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_274a_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_8dd5_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_e8f9_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_43e5_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_0215_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_6ce3_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_4430_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_a975_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_08fd_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_4dbd_return_output;
     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_060a[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_3347] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_060a_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_3347_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_060a(
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_dc8f_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_faab_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_dd63_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_8ebb_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_52da_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_87e3_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_5c81_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_a8c2_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_060a_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_3347_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
