-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity ovr_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_61914e8d;
architecture arch of ovr_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l297_c6_b407]
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l297_c2_fd37]
signal t8_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_fd37]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l297_c2_fd37]
signal n8_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l310_c11_e402]
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l310_c7_4151]
signal t8_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_4151]
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_4151]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l310_c7_4151]
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_4151]
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_4151]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l310_c7_4151]
signal n8_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l313_c11_2e62]
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l313_c7_73bc]
signal t8_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_73bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_73bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l313_c7_73bc]
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_73bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_73bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l313_c7_73bc]
signal n8_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l315_c30_f0b7]
signal sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l320_c11_d3b1]
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_c04f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_c04f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_c04f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l320_c7_c04f]
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l320_c7_c04f]
signal n8_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l326_c11_aeba]
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_c405]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_c405]
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l326_c7_c405]
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_71f0( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_left,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_right,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output);

-- t8_MUX_uxn_opcodes_h_l297_c2_fd37
t8_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
t8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
t8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37
result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- n8_MUX_uxn_opcodes_h_l297_c2_fd37
n8_MUX_uxn_opcodes_h_l297_c2_fd37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l297_c2_fd37_cond,
n8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue,
n8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse,
n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402
BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_left,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_right,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output);

-- t8_MUX_uxn_opcodes_h_l310_c7_4151
t8_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l310_c7_4151_cond,
t8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
t8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151
result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_cond,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- n8_MUX_uxn_opcodes_h_l310_c7_4151
n8_MUX_uxn_opcodes_h_l310_c7_4151 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l310_c7_4151_cond,
n8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue,
n8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse,
n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62
BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_left,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_right,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output);

-- t8_MUX_uxn_opcodes_h_l313_c7_73bc
t8_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
t8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
t8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc
result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- n8_MUX_uxn_opcodes_h_l313_c7_73bc
n8_MUX_uxn_opcodes_h_l313_c7_73bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l313_c7_73bc_cond,
n8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue,
n8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse,
n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7
sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_ins,
sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_x,
sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_y,
sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1
BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_left,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_right,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_cond,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output);

-- n8_MUX_uxn_opcodes_h_l320_c7_c04f
n8_MUX_uxn_opcodes_h_l320_c7_c04f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l320_c7_c04f_cond,
n8_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue,
n8_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse,
n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba
BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_left,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_right,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405
result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_cond,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output,
 t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output,
 t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output,
 t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output,
 sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output,
 n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_4e12 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_5df7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_3c60 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_74c2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_4019 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_e18d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_b3f7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_c405_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_4526_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_d1c5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_3572_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l332_l293_DUPLICATE_e24a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_5df7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_5df7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_b3f7 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_b3f7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_3c60 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_3c60;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_e18d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_e18d;
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_right := to_unsigned(4, 3);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_74c2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_74c2;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_4019 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_4019;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_4e12 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_4e12;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_d1c5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_d1c5_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l320_c11_d3b1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_left;
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output := BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_fd37_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l315_c30_f0b7] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_ins;
     sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_x <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_x;
     sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_y <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output := sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_fd37_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_fd37_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l313_c11_2e62] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_left;
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output := BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_4526 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_4526_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l297_c6_b407] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_left;
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output := BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l310_c11_e402] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_left;
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output := BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_fd37_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l326_c11_aeba] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_left;
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output := BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l326_c7_c405] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_c405_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_3572 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_3572_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b407_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_e402_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_2e62_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_d3b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_aeba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_3572_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_3572_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l320_l310_l326_DUPLICATE_8094_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_d1c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_d1c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_4526_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_4526_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_4526_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_fd37_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_fd37_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_fd37_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_fd37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_c405_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_f0b7_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- t8_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     t8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     t8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- n8_MUX[uxn_opcodes_h_l320_c7_c04f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l320_c7_c04f_cond <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_cond;
     n8_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue;
     n8_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output := n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_c405] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_c405] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_c04f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l326_c7_c405] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_cond;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output := result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := VAR_n8_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_c405_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_c405_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_c405_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_t8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l320_c7_c04f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output := result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;

     -- t8_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     t8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     t8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output := t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_c04f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_c04f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- n8_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     n8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     n8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_n8_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c04f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_t8_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- n8_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     n8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     n8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output := n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- t8_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     t8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     t8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_73bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_n8_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_73bc_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output := result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- n8_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     n8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     n8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_4151] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_4151_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_fd37] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l332_l293_DUPLICATE_e24a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l332_l293_DUPLICATE_e24a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_71f0(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_fd37_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_fd37_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l332_l293_DUPLICATE_e24a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l332_l293_DUPLICATE_e24a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
