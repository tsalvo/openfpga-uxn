-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity ora_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_64d180f1;
architecture arch of ora_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1007_c6_484d]
signal BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1007_c2_1d9e]
signal t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1020_c11_e8ea]
signal BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal n8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1020_c7_02d6]
signal t8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1023_c11_3cdf]
signal BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1023_c7_0589]
signal n8_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1023_c7_0589]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1023_c7_0589]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1023_c7_0589]
signal result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1023_c7_0589]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1023_c7_0589]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1023_c7_0589]
signal t8_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1026_c11_31a3]
signal BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1026_c7_832c]
signal n8_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1026_c7_832c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1026_c7_832c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1026_c7_832c]
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1026_c7_832c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1026_c7_832c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1028_c30_9229]
signal sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1031_c21_925b]
signal BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d
BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_left,
BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_right,
BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output);

-- n8_MUX_uxn_opcodes_h_l1007_c2_1d9e
n8_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e
result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- t8_MUX_uxn_opcodes_h_l1007_c2_1d9e
t8_MUX_uxn_opcodes_h_l1007_c2_1d9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond,
t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue,
t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse,
t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea
BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_left,
BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_right,
BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output);

-- n8_MUX_uxn_opcodes_h_l1020_c7_02d6
n8_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6
result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6
result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6
result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- t8_MUX_uxn_opcodes_h_l1020_c7_02d6
t8_MUX_uxn_opcodes_h_l1020_c7_02d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond,
t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue,
t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse,
t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf
BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_left,
BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_right,
BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output);

-- n8_MUX_uxn_opcodes_h_l1023_c7_0589
n8_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
n8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
n8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589
result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- t8_MUX_uxn_opcodes_h_l1023_c7_0589
t8_MUX_uxn_opcodes_h_l1023_c7_0589 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1023_c7_0589_cond,
t8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue,
t8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse,
t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_left,
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_right,
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output);

-- n8_MUX_uxn_opcodes_h_l1026_c7_832c
n8_MUX_uxn_opcodes_h_l1026_c7_832c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1026_c7_832c_cond,
n8_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue,
n8_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse,
n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1028_c30_9229
sp_relative_shift_uxn_opcodes_h_l1028_c30_9229 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_ins,
sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_x,
sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_y,
sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b
BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_left,
BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_right,
BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output,
 n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output,
 n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output,
 n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output,
 n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1012_c3_5162 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1017_c3_6141 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1021_c3_21e0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1030_c3_7014 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_84cc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_eecd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_c879_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1023_l1026_DUPLICATE_793b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1003_l1035_DUPLICATE_a57e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1012_c3_5162 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1012_c3_5162;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1030_c3_7014 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1030_c3_7014;
     VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1017_c3_6141 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1017_c3_6141;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1021_c3_21e0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1021_c3_21e0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1023_l1026_DUPLICATE_793b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1023_l1026_DUPLICATE_793b_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_c879 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_c879_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_84cc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_84cc_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_eecd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_eecd_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1007_c6_484d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1020_c11_e8ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l1028_c30_9229] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_ins;
     sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_x;
     sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output := sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1031_c21_925b] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_left;
     BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output := BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1026_c11_31a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1023_c11_3cdf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_left;
     BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output := BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output := result.is_ram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c6_484d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1020_c11_e8ea_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c11_3cdf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_31a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1031_c21_925b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_eecd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_eecd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_eecd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_84cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_84cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_84cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_c879_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_c879_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1023_l1020_l1026_DUPLICATE_c879_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1023_l1026_DUPLICATE_793b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1023_l1026_DUPLICATE_793b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1023_l1007_l1020_l1026_DUPLICATE_f990_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1007_c2_1d9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1028_c30_9229_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1026_c7_832c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     t8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     t8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1026_c7_832c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1026_c7_832c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1026_c7_832c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1026_c7_832c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_cond;
     n8_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue;
     n8_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output := n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1026_c7_832c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1026_c7_832c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_832c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- t8_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l1023_c7_0589] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1023_c7_0589_cond <= VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_cond;
     n8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_iftrue;
     n8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output := n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1023_c7_0589_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1020_c7_02d6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;

     -- t8_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1020_c7_02d6_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1007_c2_1d9e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1003_l1035_DUPLICATE_a57e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1003_l1035_DUPLICATE_a57e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1007_c2_1d9e_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1003_l1035_DUPLICATE_a57e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1003_l1035_DUPLICATE_a57e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
