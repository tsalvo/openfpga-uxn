-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc2_0CLK_180c5210 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_180c5210;
architecture arch of inc2_0CLK_180c5210 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_463f]
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1355_c2_d559]
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1355_c2_d559]
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_d559]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_ef6a]
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1368_c7_084d]
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1368_c7_084d]
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_084d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_084d]
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_084d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_084d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_084d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_46ce]
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_eaf0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_d59a]
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output : unsigned(8 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1373_c30_64bb]
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_ff13]
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1378_c7_f13d]
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_f13d]
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_f13d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_f13d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_f13d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_b359]
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1379_c37_af46]
signal MUX_uxn_opcodes_h_l1379_c37_af46_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_af46_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_af46_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_af46_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_8da7]
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_left,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_right,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1355_c2_d559
t16_low_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1355_c2_d559
t16_high_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_left,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_right,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1368_c7_084d
t16_low_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1368_c7_084d
t16_high_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_left,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_right,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0
t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0
t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_left,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_right,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb
sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_ins,
sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_x,
sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_y,
sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_left,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_right,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d
t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_cond,
t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue,
t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse,
t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_left,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_right,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output);

-- MUX_uxn_opcodes_h_l1379_c37_af46
MUX_uxn_opcodes_h_l1379_c37_af46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1379_c37_af46_cond,
MUX_uxn_opcodes_h_l1379_c37_af46_iftrue,
MUX_uxn_opcodes_h_l1379_c37_af46_iffalse,
MUX_uxn_opcodes_h_l1379_c37_af46_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_left,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_right,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output,
 t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output,
 t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output,
 t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output,
 sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output,
 t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output,
 MUX_uxn_opcodes_h_l1379_c37_af46_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_087b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_ca91 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_7a8f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_uxn_opcodes_h_l1372_c3_92b5 : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_c831 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output : unsigned(8 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_uxn_opcodes_h_l1379_c3_df61 : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_5c84 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_457b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_f13d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_left : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_af46_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_af46_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_af46_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_af46_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_5e1b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_144d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_f13b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_fbdc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1386_l1351_DUPLICATE_d6b3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_5c84 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_5c84;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_ca91 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_ca91;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1379_c37_af46_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_7a8f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_7a8f;
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_MUX_uxn_opcodes_h_l1379_c37_af46_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_right := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_457b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_457b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_c831 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_c831;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_087b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_087b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_left := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_left := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse := t16_high;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_left := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := t16_low;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_d559_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_5e1b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_5e1b_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1378_c7_f13d] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_f13d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_b359] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_left;
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output := BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_144d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_144d_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_d559_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_46ce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_left;
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output := BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_ff13] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_left;
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output := BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_f13b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_f13b_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_d559_return_output := result.is_ram_write;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_d59a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_ef6a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_d559_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_fbdc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_fbdc_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1373_c30_64bb] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_ins;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_x;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output := sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_463f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_463f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_ef6a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_46ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_ff13_return_output;
     VAR_MUX_uxn_opcodes_h_l1379_c37_af46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_b359_return_output;
     VAR_t16_low_uxn_opcodes_h_l1372_c3_92b5 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_d59a_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_f13b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_f13b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_fbdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_fbdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_fbdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_144d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_144d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_5e1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_5e1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_5e1b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_d559_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_d559_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_d559_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_d559_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_f13d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_64bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_92b5;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_92b5;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_f13d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_f13d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;

     -- MUX[uxn_opcodes_h_l1379_c37_af46] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1379_c37_af46_cond <= VAR_MUX_uxn_opcodes_h_l1379_c37_af46_cond;
     MUX_uxn_opcodes_h_l1379_c37_af46_iftrue <= VAR_MUX_uxn_opcodes_h_l1379_c37_af46_iftrue;
     MUX_uxn_opcodes_h_l1379_c37_af46_iffalse <= VAR_MUX_uxn_opcodes_h_l1379_c37_af46_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1379_c37_af46_return_output := MUX_uxn_opcodes_h_l1379_c37_af46_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_f13d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_right := VAR_MUX_uxn_opcodes_h_l1379_c37_af46_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_8da7] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output;

     -- Submodule level 3
     VAR_t16_high_uxn_opcodes_h_l1379_c3_df61 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_8da7_return_output, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_df61;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_df61;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_f13d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1378_c7_f13d] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_cond;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output := t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_f13d_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1371_c7_eaf0] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_cond;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output := t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_eaf0_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_084d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_084d_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_d559] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output := result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;

     -- Submodule level 7
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_d559_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1386_l1351_DUPLICATE_d6b3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1386_l1351_DUPLICATE_d6b3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_d559_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_d559_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1386_l1351_DUPLICATE_d6b3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1386_l1351_DUPLICATE_d6b3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
