-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity and_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_64d180f1;
architecture arch of and_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l927_c6_f5ad]
signal BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l927_c2_8c76]
signal t8_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l927_c2_8c76]
signal n8_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l927_c2_8c76]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l940_c11_dd9c]
signal BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l940_c7_b99c]
signal t8_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l940_c7_b99c]
signal n8_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l940_c7_b99c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l940_c7_b99c]
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l940_c7_b99c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l940_c7_b99c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l940_c7_b99c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l943_c11_bf19]
signal BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l943_c7_19fb]
signal t8_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l943_c7_19fb]
signal n8_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l943_c7_19fb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l943_c7_19fb]
signal result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l943_c7_19fb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l943_c7_19fb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l943_c7_19fb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l946_c11_0523]
signal BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l946_c7_b625]
signal n8_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l946_c7_b625]
signal result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l946_c7_b625]
signal result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l946_c7_b625]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l946_c7_b625]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l946_c7_b625]
signal result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l948_c30_bdc7]
signal sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l951_c21_fa38]
signal BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad
BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_left,
BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_right,
BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output);

-- t8_MUX_uxn_opcodes_h_l927_c2_8c76
t8_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
t8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
t8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- n8_MUX_uxn_opcodes_h_l927_c2_8c76
n8_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
n8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
n8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76
result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76
result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76
result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76
result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76
result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76
result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76
result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c
BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_left,
BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_right,
BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output);

-- t8_MUX_uxn_opcodes_h_l940_c7_b99c
t8_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
t8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
t8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- n8_MUX_uxn_opcodes_h_l940_c7_b99c
n8_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
n8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
n8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c
result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19
BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_left,
BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_right,
BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output);

-- t8_MUX_uxn_opcodes_h_l943_c7_19fb
t8_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
t8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
t8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- n8_MUX_uxn_opcodes_h_l943_c7_19fb
n8_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
n8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
n8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb
result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb
result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb
result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb
result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523
BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_left,
BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_right,
BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output);

-- n8_MUX_uxn_opcodes_h_l946_c7_b625
n8_MUX_uxn_opcodes_h_l946_c7_b625 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l946_c7_b625_cond,
n8_MUX_uxn_opcodes_h_l946_c7_b625_iftrue,
n8_MUX_uxn_opcodes_h_l946_c7_b625_iffalse,
n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625
result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625
result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_cond,
result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625
result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625
result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output);

-- sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7
sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_ins,
sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_x,
sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_y,
sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38
BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_left,
BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_right,
BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output,
 t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output,
 t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output,
 t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output,
 n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output,
 sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output,
 BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l932_c3_54fd : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l937_c3_b617 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l941_c3_ad1f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l950_c3_4e35 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_81b9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_6ada_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_3863_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l943_l946_DUPLICATE_1e48_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l955_l923_DUPLICATE_b11d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l950_c3_4e35 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l950_c3_4e35;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l932_c3_54fd := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l932_c3_54fd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l941_c3_ad1f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l941_c3_ad1f;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l937_c3_b617 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l937_c3_b617;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := t8;
     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l927_c2_8c76_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l927_c2_8c76_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l943_l946_DUPLICATE_1e48 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l943_l946_DUPLICATE_1e48_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l927_c2_8c76_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l927_c6_f5ad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_left;
     BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output := BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_81b9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_81b9_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_6ada LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_6ada_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l948_c30_bdc7] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_ins;
     sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_x <= VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_x;
     sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_y <= VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output := sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l940_c11_dd9c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_left;
     BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output := BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l927_c2_8c76_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l943_c11_bf19] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_left;
     BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output := BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l946_c11_0523] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_left;
     BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output := BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l951_c21_fa38] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_left;
     BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output := BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_3863 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_3863_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l951_c21_fa38_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l927_c6_f5ad_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_dd9c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l943_c11_bf19_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l946_c11_0523_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_6ada_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_6ada_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_6ada_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_81b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_81b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_81b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_3863_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_3863_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l943_l946_l940_DUPLICATE_3863_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l943_l946_DUPLICATE_1e48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l943_l946_DUPLICATE_1e48_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l943_l946_l940_l927_DUPLICATE_f22d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l927_c2_8c76_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l927_c2_8c76_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l927_c2_8c76_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l927_c2_8c76_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l948_c30_bdc7_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l946_c7_b625] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l946_c7_b625] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l946_c7_b625] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l946_c7_b625] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_cond;
     result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output := result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- n8_MUX[uxn_opcodes_h_l946_c7_b625] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l946_c7_b625_cond <= VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_cond;
     n8_MUX_uxn_opcodes_h_l946_c7_b625_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_iftrue;
     n8_MUX_uxn_opcodes_h_l946_c7_b625_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output := n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l946_c7_b625] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output;

     -- t8_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     t8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     t8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l946_c7_b625_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l946_c7_b625_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l946_c7_b625_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l946_c7_b625_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l946_c7_b625_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l946_c7_b625_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     -- n8_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     n8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     n8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- t8_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     t8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     t8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l943_c7_19fb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l943_c7_19fb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_t8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     -- t8_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     t8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     t8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- n8_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     n8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     n8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l940_c7_b99c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_n8_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_b99c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- n8_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     n8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     n8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l927_c2_8c76] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l927_c2_8c76_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l955_l923_DUPLICATE_b11d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l955_l923_DUPLICATE_b11d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l927_c2_8c76_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l927_c2_8c76_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l955_l923_DUPLICATE_b11d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l955_l923_DUPLICATE_b11d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
