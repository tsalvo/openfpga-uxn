-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity ora_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_bacf6a1d;
architecture arch of ora_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l956_c6_52d7]
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_9fac]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l956_c2_741e]
signal n8_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l956_c2_741e]
signal t8_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_741e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_741e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_741e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_741e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_741e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l956_c2_741e]
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l957_c3_56f0[uxn_opcodes_h_l957_c3_56f0]
signal printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l961_c11_41c0]
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal n8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal t8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l961_c7_c4e0]
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l964_c11_b85c]
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal n8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal t8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l964_c7_e7c8]
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l967_c11_c1d6]
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal n8_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l967_c7_6ee9]
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l970_c30_677f]
signal sp_relative_shift_uxn_opcodes_h_l970_c30_677f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_677f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_677f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l973_c21_a361]
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l975_c11_92d9]
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_575d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_575d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_575d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7
BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_left,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_right,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output);

-- n8_MUX_uxn_opcodes_h_l956_c2_741e
n8_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l956_c2_741e_cond,
n8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
n8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- t8_MUX_uxn_opcodes_h_l956_c2_741e
t8_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l956_c2_741e_cond,
t8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
t8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e
result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_cond,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

-- printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0
printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0 : entity work.printf_uxn_opcodes_h_l957_c3_56f0_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0
BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_left,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_right,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output);

-- n8_MUX_uxn_opcodes_h_l961_c7_c4e0
n8_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- t8_MUX_uxn_opcodes_h_l961_c7_c4e0
t8_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_cond,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c
BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_left,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_right,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output);

-- n8_MUX_uxn_opcodes_h_l964_c7_e7c8
n8_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- t8_MUX_uxn_opcodes_h_l964_c7_e7c8
t8_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8
result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_cond,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6
BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_left,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_right,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output);

-- n8_MUX_uxn_opcodes_h_l967_c7_6ee9
n8_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9
result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_cond,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l970_c30_677f
sp_relative_shift_uxn_opcodes_h_l970_c30_677f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l970_c30_677f_ins,
sp_relative_shift_uxn_opcodes_h_l970_c30_677f_x,
sp_relative_shift_uxn_opcodes_h_l970_c30_677f_y,
sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l973_c21_a361
BIN_OP_OR_uxn_opcodes_h_l973_c21_a361 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_left,
BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_right,
BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9
BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_left,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_right,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output,
 n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output,
 n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output,
 n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output,
 n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output,
 sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output,
 BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_b6b3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_d817 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_d922 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_4b89_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l981_l952_DUPLICATE_dd4a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_b6b3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_b6b3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_d817 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_d817;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_d922 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_d922;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_y := resize(to_signed(-1, 2), 4);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l967_c11_c1d6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_left;
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output := BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l961_c11_41c0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_left;
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output := BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l964_c11_b85c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_left;
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output := BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l956_c6_52d7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_left;
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output := BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l970_c30_677f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l970_c30_677f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_ins;
     sp_relative_shift_uxn_opcodes_h_l970_c30_677f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_x;
     sp_relative_shift_uxn_opcodes_h_l970_c30_677f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output := sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l975_c11_92d9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_left;
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output := BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1_return_output := result.is_stack_write;

     -- BIN_OP_OR[uxn_opcodes_h_l973_c21_a361] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_left;
     BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output := BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_4b89 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_4b89_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_52d7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_41c0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_b85c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_c1d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_92d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_a361_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_b24a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l975_l964_l967_l961_DUPLICATE_af5a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_41bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l975_l964_l956_l961_DUPLICATE_9db1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_4b89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_4b89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_195d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_677f_return_output;
     -- n8_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_9fac] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_575d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_575d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output;

     -- t8_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_575d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_9fac_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_575d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_575d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_575d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     -- n8_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- printf_uxn_opcodes_h_l957_c3_56f0[uxn_opcodes_h_l957_c3_56f0] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l957_c3_56f0_uxn_opcodes_h_l957_c3_56f0_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- t8_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_6ee9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_6ee9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- n8_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_e7c8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;

     -- t8_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     t8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     t8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output := t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_e7c8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l956_c2_741e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output := result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- n8_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     n8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     n8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output := n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_c4e0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l956_c2_741e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c4e0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_741e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l981_l952_DUPLICATE_dd4a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l981_l952_DUPLICATE_dd4a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_741e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_741e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l981_l952_DUPLICATE_dd4a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l981_l952_DUPLICATE_dd4a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
