-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity mul2_0CLK_06b39b76 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end mul2_0CLK_06b39b76;
architecture arch of mul2_0CLK_06b39b76 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1826_c6_4e25]
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal n16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1826_c2_b15a]
signal t16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1834_c11_1bda]
signal BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1834_c7_2871]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1834_c7_2871]
signal n16_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1834_c7_2871]
signal tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1834_c7_2871]
signal t16_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1837_c11_d06f]
signal BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal n16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1837_c7_57ec]
signal t16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1840_c30_0d5c]
signal sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1842_c11_cae4]
signal BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal n16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1842_c7_08a1]
signal tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(15 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1844_c11_9e15]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_left : unsigned(15 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_right : unsigned(15 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1850_c11_7822]
signal BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1850_c7_1985]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1850_c7_1985]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1850_c7_1985]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_left,
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_right,
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a
result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a
result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- n16_MUX_uxn_opcodes_h_l1826_c2_b15a
n16_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a
tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- t16_MUX_uxn_opcodes_h_l1826_c2_b15a
t16_MUX_uxn_opcodes_h_l1826_c2_b15a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond,
t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue,
t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse,
t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda
BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_left,
BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_right,
BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871
result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871
result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871
result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871
result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871
result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- n16_MUX_uxn_opcodes_h_l1834_c7_2871
n16_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
n16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
n16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1834_c7_2871
tmp16_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- t16_MUX_uxn_opcodes_h_l1834_c7_2871
t16_MUX_uxn_opcodes_h_l1834_c7_2871 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1834_c7_2871_cond,
t16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue,
t16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse,
t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f
BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_left,
BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_right,
BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec
result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec
result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec
result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec
result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec
result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- n16_MUX_uxn_opcodes_h_l1837_c7_57ec
n16_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec
tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- t16_MUX_uxn_opcodes_h_l1837_c7_57ec
t16_MUX_uxn_opcodes_h_l1837_c7_57ec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond,
t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue,
t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse,
t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c
sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_ins,
sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_x,
sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_y,
sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_left,
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_right,
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1
result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1
result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- n16_MUX_uxn_opcodes_h_l1842_c7_08a1
n16_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1
tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond,
tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue,
tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse,
tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15 : entity work.BIN_OP_INFERRED_MULT_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822
BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_left,
BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_right,
BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985
result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985
result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output,
 sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1831_c3_787a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1835_c3_9e31 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1847_c3_3b81 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_uxn_opcodes_h_l1844_c3_0269 : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1842_l1834_l1826_DUPLICATE_5ef8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1834_l1837_l1826_DUPLICATE_e857_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1837_DUPLICATE_d74e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1856_l1822_DUPLICATE_1730_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1835_c3_9e31 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1835_c3_9e31;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1831_c3_787a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1831_c3_787a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_right := to_unsigned(4, 3);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1847_c3_3b81 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1847_c3_3b81;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := t16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l1837_c11_d06f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1834_l1837_l1826_DUPLICATE_e857 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1834_l1837_l1826_DUPLICATE_e857_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1834_c11_1bda] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_left;
     BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output := BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1826_c6_4e25] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_left;
     BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output := BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1842_l1834_l1826_DUPLICATE_5ef8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1842_l1834_l1826_DUPLICATE_5ef8_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1840_c30_0d5c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_ins;
     sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_x;
     sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output := sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1850_c11_7822] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_left;
     BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output := BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1844_c11_9e15] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1842_c11_cae4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1837_DUPLICATE_d74e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1837_DUPLICATE_d74e_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_4e25_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1834_c11_1bda_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1837_c11_d06f_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_cae4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1850_c11_7822_return_output;
     VAR_tmp16_uxn_opcodes_h_l1844_c3_0269 := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1844_c11_9e15_return_output, 16);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1834_l1837_l1826_DUPLICATE_e857_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1834_l1837_l1826_DUPLICATE_e857_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1834_l1837_l1826_DUPLICATE_e857_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1842_l1834_l1837_l1826_DUPLICATE_a619_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_c7a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1842_l1834_l1826_DUPLICATE_5ef8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1842_l1834_l1826_DUPLICATE_5ef8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1842_l1834_l1826_DUPLICATE_5ef8_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1842_l1834_l1850_l1837_DUPLICATE_8a0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1834_l1850_l1837_l1826_DUPLICATE_c8be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1837_DUPLICATE_d74e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1837_DUPLICATE_d74e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1840_c30_0d5c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := VAR_tmp16_uxn_opcodes_h_l1844_c3_0269;
     VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue := VAR_tmp16_uxn_opcodes_h_l1844_c3_0269;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1850_c7_1985] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- n16_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1850_c7_1985] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1850_c7_1985] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output;

     -- t16_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1850_c7_1985_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1850_c7_1985_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1850_c7_1985_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- t16_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     t16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     t16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1842_c7_08a1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- n16_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_08a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- n16_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     n16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     n16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- t16_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1837_c7_57ec] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1837_c7_57ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1834_c7_2871] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;

     -- n16_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1834_c7_2871_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1826_c2_b15a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1856_l1822_DUPLICATE_1730 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1856_l1822_DUPLICATE_1730_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_b15a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1856_l1822_DUPLICATE_1730_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1856_l1822_DUPLICATE_1730_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
