-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity gth_0CLK_57104a4d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_57104a4d;
architecture arch of gth_0CLK_57104a4d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1919_c6_8da5]
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1919_c2_1eb4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1924_c11_d051]
signal BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal n8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal t8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1924_c7_5e35]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1927_c11_faa7]
signal BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1927_c7_0174]
signal n8_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1927_c7_0174]
signal t8_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1927_c7_0174]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1927_c7_0174]
signal result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1927_c7_0174]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1927_c7_0174]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1927_c7_0174]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1927_c7_0174]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_a488]
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1931_c7_d2ef]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1934_c11_da8f]
signal BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal n8_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1934_c7_8e57]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1937_c30_9e4d]
signal sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1940_c21_bd4e]
signal BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1940_c21_956b]
signal MUX_uxn_opcodes_h_l1940_c21_956b_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1940_c21_956b_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1940_c21_956b_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1940_c21_956b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1942_c11_215e]
signal BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1942_c7_9e0b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1942_c7_9e0b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1942_c7_9e0b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5
BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_left,
BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_right,
BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output);

-- n8_MUX_uxn_opcodes_h_l1919_c2_1eb4
n8_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- t8_MUX_uxn_opcodes_h_l1919_c2_1eb4
t8_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4
result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4
result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_left,
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_right,
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output);

-- n8_MUX_uxn_opcodes_h_l1924_c7_5e35
n8_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- t8_MUX_uxn_opcodes_h_l1924_c7_5e35
t8_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7
BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_left,
BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_right,
BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output);

-- n8_MUX_uxn_opcodes_h_l1927_c7_0174
n8_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
n8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
n8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- t8_MUX_uxn_opcodes_h_l1927_c7_0174
t8_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
t8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
t8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174
result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174
result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174
result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174
result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174
result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_left,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_right,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output);

-- n8_MUX_uxn_opcodes_h_l1931_c7_d2ef
n8_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f
BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_left,
BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_right,
BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output);

-- n8_MUX_uxn_opcodes_h_l1934_c7_8e57
n8_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57
result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57
result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57
result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57
result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57
result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d
sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_ins,
sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_x,
sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_y,
sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e
BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_left,
BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_right,
BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output);

-- MUX_uxn_opcodes_h_l1940_c21_956b
MUX_uxn_opcodes_h_l1940_c21_956b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1940_c21_956b_cond,
MUX_uxn_opcodes_h_l1940_c21_956b_iftrue,
MUX_uxn_opcodes_h_l1940_c21_956b_iffalse,
MUX_uxn_opcodes_h_l1940_c21_956b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e
BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_left,
BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_right,
BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b
result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b
result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b
result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output,
 n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output,
 n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output,
 n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output,
 n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output,
 n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output,
 sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output,
 MUX_uxn_opcodes_h_l1940_c21_956b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1921_c3_5fc0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1925_c3_295d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_e5fa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1932_c3_65bf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1939_c3_6624 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1934_c7_8e57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1940_c21_956b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1940_c21_956b_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1940_c21_956b_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1940_c21_956b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1948_l1915_DUPLICATE_cc23_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1921_c3_5fc0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1921_c3_5fc0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_e5fa := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_e5fa;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1940_c21_956b_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1932_c3_65bf := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1932_c3_65bf;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1940_c21_956b_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1939_c3_6624 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1939_c3_6624;
     VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1925_c3_295d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1925_c3_295d;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_a488] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_left;
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output := BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1942_c11_215e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1927_c11_faa7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1924_c11_d051] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_left;
     BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output := BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1919_c6_8da5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1934_c11_da8f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output := result.sp_relative_shift;

     -- BIN_OP_GT[uxn_opcodes_h_l1940_c21_bd4e] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_left;
     BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output := BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1934_c7_8e57_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1937_c30_9e4d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_ins;
     sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_x;
     sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output := sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c6_8da5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_d051_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1927_c11_faa7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_a488_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1934_c11_da8f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1942_c11_215e_return_output;
     VAR_MUX_uxn_opcodes_h_l1940_c21_956b_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1940_c21_bd4e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_d15d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1942_l1934_DUPLICATE_bcb2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_1e7d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1942_DUPLICATE_18a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1931_l1927_l1924_l1919_l1934_DUPLICATE_a91e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1937_c30_9e4d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- n8_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1942_c7_9e0b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1942_c7_9e0b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1942_c7_9e0b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output;

     -- MUX[uxn_opcodes_h_l1940_c21_956b] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1940_c21_956b_cond <= VAR_MUX_uxn_opcodes_h_l1940_c21_956b_cond;
     MUX_uxn_opcodes_h_l1940_c21_956b_iftrue <= VAR_MUX_uxn_opcodes_h_l1940_c21_956b_iftrue;
     MUX_uxn_opcodes_h_l1940_c21_956b_iffalse <= VAR_MUX_uxn_opcodes_h_l1940_c21_956b_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1940_c21_956b_return_output := MUX_uxn_opcodes_h_l1940_c21_956b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     t8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     t8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue := VAR_MUX_uxn_opcodes_h_l1940_c21_956b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1942_c7_9e0b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- n8_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- t8_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1934_c7_8e57] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1934_c7_8e57_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     -- n8_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     n8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     n8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- t8_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1931_c7_d2ef] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_d2ef_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- n8_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1927_c7_0174] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1927_c7_0174_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1924_c7_5e35] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_5e35_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1919_c2_1eb4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1948_l1915_DUPLICATE_cc23 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1948_l1915_DUPLICATE_cc23_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1919_c2_1eb4_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1948_l1915_DUPLICATE_cc23_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1948_l1915_DUPLICATE_cc23_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
