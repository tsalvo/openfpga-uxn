-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ldr_0CLK_46731a7b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_46731a7b;
architecture arch of ldr_0CLK_46731a7b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1692_c6_f98f]
signal BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal t8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1692_c2_22d0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1697_c11_6b7f]
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal t8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1697_c7_14f0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1700_c11_8c7f]
signal BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1700_c7_1826]
signal tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1700_c7_1826]
signal t8_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1700_c7_1826]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1703_c30_2068]
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1704_c22_e9cf]
signal BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1706_c11_6479]
signal BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1706_c7_30c6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1708_c22_d44a]
signal BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1710_c11_1a09]
signal BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1710_c7_9217]
signal tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1710_c7_9217]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1710_c7_9217]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1710_c7_9217]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1710_c7_9217]
signal result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1716_c11_7a5f]
signal BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1716_c7_d277]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1716_c7_d277]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_sp_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f
BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_left,
BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_right,
BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0
tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- t8_MUX_uxn_opcodes_h_l1692_c2_22d0
t8_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0
result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0
result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0
result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0
result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0
result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_left,
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_right,
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0
tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- t8_MUX_uxn_opcodes_h_l1697_c7_14f0
t8_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_left,
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_right,
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1700_c7_1826
tmp8_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- t8_MUX_uxn_opcodes_h_l1700_c7_1826
t8_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
t8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
t8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826
result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826
result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1703_c30_2068
sp_relative_shift_uxn_opcodes_h_l1703_c30_2068 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_ins,
sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_x,
sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_y,
sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf
BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_left,
BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_right,
BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_left,
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_right,
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6
tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6
result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6
result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a
BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_left,
BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_right,
BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09
BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_left,
BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_right,
BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1710_c7_9217
tmp8_MUX_uxn_opcodes_h_l1710_c7_9217 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_cond,
tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue,
tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse,
tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217
result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217
result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217
result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_cond,
result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f
BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_left,
BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_right,
BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277
result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277
result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output,
 sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output,
 tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output,
 tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1694_c3_d577 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1698_c3_26d2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1704_c3_ee34 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1704_c27_d101_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1708_c3_5659 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1708_c27_3333_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1713_c3_827c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_491b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1692_l1697_l1700_DUPLICATE_868f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_3062_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1706_l1710_l1700_DUPLICATE_b330_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1721_l1688_DUPLICATE_4477_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1713_c3_827c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1713_c3_827c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1694_c3_d577 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1694_c3_d577;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1698_c3_26d2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1698_c3_26d2;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1697_c11_6b7f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1703_c30_2068] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_ins;
     sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_x;
     sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output := sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1692_c6_f98f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_3062 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_3062_return_output := result.is_sp_shift;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1708_c27_3333] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1708_c27_3333_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1706_c11_6479] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_left;
     BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output := BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1692_l1697_l1700_DUPLICATE_868f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1692_l1697_l1700_DUPLICATE_868f_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1716_c11_7a5f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_491b LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_491b_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1700_c11_8c7f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1710_c11_1a09] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_left;
     BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output := BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1704_c27_d101] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1704_c27_d101_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1706_l1710_l1700_DUPLICATE_b330 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1706_l1710_l1700_DUPLICATE_b330_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1692_c6_f98f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_6b7f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_8c7f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6479_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1710_c11_1a09_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1716_c11_7a5f_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1704_c27_d101_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1708_c27_3333_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1692_l1697_l1700_DUPLICATE_868f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1692_l1697_l1700_DUPLICATE_868f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1692_l1697_l1700_DUPLICATE_868f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_491b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_491b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_491b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1716_l1710_l1706_l1700_l1697_DUPLICATE_20b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_3062_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_3062_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1692_l1706_l1697_DUPLICATE_3062_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1692_l1716_l1706_l1700_l1697_DUPLICATE_e83a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1706_l1710_l1700_DUPLICATE_b330_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1706_l1710_l1700_DUPLICATE_b330_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1706_l1710_l1700_DUPLICATE_b330_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1692_l1710_l1706_l1700_l1697_DUPLICATE_51dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_2068_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1716_c7_d277] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1704_c22_e9cf] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1710_c7_9217] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;

     -- t8_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     t8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     t8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1716_c7_d277] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1708_c22_d44a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1710_c7_9217] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_cond;
     tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output := tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1710_c7_9217] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output := result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1704_c3_ee34 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1704_c22_e9cf_return_output)),16);
     VAR_result_u16_value_uxn_opcodes_h_l1708_c3_5659 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1708_c22_d44a_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1716_c7_d277_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1716_c7_d277_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1704_c3_ee34;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1708_c3_5659;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1710_c7_9217] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;

     -- t8_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1710_c7_9217] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1710_c7_9217_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1706_c7_30c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1706_c7_30c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1700_c7_1826] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1700_c7_1826_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1697_c7_14f0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_14f0_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1692_c2_22d0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1721_l1688_DUPLICATE_4477 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1721_l1688_DUPLICATE_4477_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1692_c2_22d0_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1721_l1688_DUPLICATE_4477_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1721_l1688_DUPLICATE_4477_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
