-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity opc_ldr_phased_0CLK_0753a953 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_ldr_phased_0CLK_0753a953;
architecture arch of opc_ldr_phased_0CLK_0753a953 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal ram8_at_tmp16 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp16 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_t8 : unsigned(15 downto 0);
signal REG_COMB_ram8_at_tmp16 : unsigned(7 downto 0);
signal REG_COMB_tmp16 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l742_c6_f79e]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l742_c1_d064]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l745_c7_65a3]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l742_c2_e567]
signal t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(15 downto 0);

-- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l742_c2_e567]
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_phased_h_l742_c2_e567]
signal tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(7 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(7 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l742_c2_e567]
signal result_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l743_c12_200c]
signal set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l745_c11_cd5f]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l745_c1_9e5b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l748_c7_2112]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l745_c7_65a3]
signal t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(15 downto 0);

-- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l745_c7_65a3]
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_phased_h_l745_c7_65a3]
signal tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(7 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(7 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l745_c7_65a3]
signal result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l746_c8_d4e1]
signal t_register_uxn_opcodes_phased_h_l746_c8_d4e1_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l748_c11_364d]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l748_c1_72a3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l753_c7_28d0]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l748_c7_2112]
signal t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(15 downto 0);

-- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l748_c7_2112]
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_phased_h_l748_c7_2112]
signal tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(7 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(7 downto 0);
signal tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l748_c7_2112]
signal result_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l749_c8_5b93]
signal t_register_uxn_opcodes_phased_h_l749_c8_5b93_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_phased_h_l750_c11_aeb5]
signal BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output : signed(17 downto 0);

-- peek_ram[uxn_opcodes_phased_h_l751_c19_a4da]
signal peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_CLOCK_ENABLE : unsigned(0 downto 0);
signal peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_address : unsigned(15 downto 0);
signal peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l753_c11_24df]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l753_c1_1c15]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l757_c7_5795]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output : unsigned(0 downto 0);

-- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l753_c7_28d0]
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond : unsigned(0 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse : unsigned(7 downto 0);
signal ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l753_c7_28d0]
signal result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output : unsigned(0 downto 0);

-- peek_ram[uxn_opcodes_phased_h_l754_c19_6dee]
signal peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_CLOCK_ENABLE : unsigned(0 downto 0);
signal peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_address : unsigned(15 downto 0);
signal peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output : unsigned(7 downto 0);

-- set[uxn_opcodes_phased_h_l755_c3_0b69]
signal set_uxn_opcodes_phased_h_l755_c3_0b69_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l755_c3_0b69_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l755_c3_0b69_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l755_c3_0b69_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l755_c3_0b69_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l755_c3_0b69_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l755_c3_0b69_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l757_c11_cef8]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l757_c1_0057]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l757_c7_5795]
signal result_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_phased_h_l758_c3_d8d5]
signal put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l760_c11_169d]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l760_c7_9071]
signal result_MUX_uxn_opcodes_phased_h_l760_c7_9071_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint16_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e
BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l742_c2_e567
t8_MUX_uxn_opcodes_phased_h_l742_c2_e567 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond,
t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue,
t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse,
t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output);

-- ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output);

-- tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567
tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond,
tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue,
tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse,
tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output);

-- result_MUX_uxn_opcodes_phased_h_l742_c2_e567
result_MUX_uxn_opcodes_phased_h_l742_c2_e567 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond,
result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue,
result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse,
result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l743_c12_200c
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_sp,
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_k,
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_mul,
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_add,
set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f
BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3
t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond,
t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue,
t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse,
t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output);

-- ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output);

-- tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3
tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond,
tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue,
tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse,
tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output);

-- result_MUX_uxn_opcodes_phased_h_l745_c7_65a3
result_MUX_uxn_opcodes_phased_h_l745_c7_65a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond,
result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue,
result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse,
result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output);

-- t_register_uxn_opcodes_phased_h_l746_c8_d4e1
t_register_uxn_opcodes_phased_h_l746_c8_d4e1 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l746_c8_d4e1_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_index,
t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_ptr,
t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d
BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l748_c7_2112
t8_MUX_uxn_opcodes_phased_h_l748_c7_2112 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond,
t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue,
t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse,
t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output);

-- ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output);

-- tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112
tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond,
tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue,
tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse,
tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output);

-- result_MUX_uxn_opcodes_phased_h_l748_c7_2112
result_MUX_uxn_opcodes_phased_h_l748_c7_2112 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond,
result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue,
result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse,
result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output);

-- t_register_uxn_opcodes_phased_h_l749_c8_5b93
t_register_uxn_opcodes_phased_h_l749_c8_5b93 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l749_c8_5b93_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_index,
t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_ptr,
t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output);

-- BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5
BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_left,
BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_right,
BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output);

-- peek_ram_uxn_opcodes_phased_h_l751_c19_a4da
peek_ram_uxn_opcodes_phased_h_l751_c19_a4da : entity work.peek_ram_0CLK_7bf2eff3 port map (
clk,
peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_CLOCK_ENABLE,
peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_address,
peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df
BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output);

-- ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse,
ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output);

-- result_MUX_uxn_opcodes_phased_h_l753_c7_28d0
result_MUX_uxn_opcodes_phased_h_l753_c7_28d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond,
result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue,
result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse,
result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output);

-- peek_ram_uxn_opcodes_phased_h_l754_c19_6dee
peek_ram_uxn_opcodes_phased_h_l754_c19_6dee : entity work.peek_ram_0CLK_7bf2eff3 port map (
clk,
peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_CLOCK_ENABLE,
peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_address,
peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output);

-- set_uxn_opcodes_phased_h_l755_c3_0b69
set_uxn_opcodes_phased_h_l755_c3_0b69 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l755_c3_0b69_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l755_c3_0b69_sp,
set_uxn_opcodes_phased_h_l755_c3_0b69_stack_index,
set_uxn_opcodes_phased_h_l755_c3_0b69_ins,
set_uxn_opcodes_phased_h_l755_c3_0b69_k,
set_uxn_opcodes_phased_h_l755_c3_0b69_mul,
set_uxn_opcodes_phased_h_l755_c3_0b69_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8
BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output);

-- result_MUX_uxn_opcodes_phased_h_l757_c7_5795
result_MUX_uxn_opcodes_phased_h_l757_c7_5795 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond,
result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue,
result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse,
result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output);

-- put_stack_uxn_opcodes_phased_h_l758_c3_d8d5
put_stack_uxn_opcodes_phased_h_l758_c3_d8d5 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_sp,
put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_stack_index,
put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_offset,
put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d
BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output);

-- result_MUX_uxn_opcodes_phased_h_l760_c7_9071
result_MUX_uxn_opcodes_phased_h_l760_c7_9071 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l760_c7_9071_cond,
result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iftrue,
result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iffalse,
result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 t8,
 ram8_at_tmp16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output,
 t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output,
 ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output,
 tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output,
 result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output,
 set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output,
 t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output,
 ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output,
 tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output,
 result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output,
 t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output,
 t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output,
 ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output,
 tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output,
 result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output,
 t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output,
 BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output,
 peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output,
 ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output,
 result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output,
 peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output,
 result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output,
 result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(15 downto 0);
 variable VAR_t8_uxn_opcodes_phased_h_l746_c3_f1e4 : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(15 downto 0);
 variable VAR_t8_uxn_opcodes_phased_h_l749_c3_4ab4 : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(7 downto 0);
 variable VAR_tmp16_uxn_opcodes_phased_h_l750_c3_ceda : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(7 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_phased_h_l750_c17_1f12_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output : signed(17 downto 0);
 variable VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_address : unsigned(15 downto 0);
 variable VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse : unsigned(0 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse : unsigned(7 downto 0);
 variable VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond : unsigned(0 downto 0);
 variable VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_address : unsigned(15 downto 0);
 variable VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(15 downto 0);
variable REG_VAR_ram8_at_tmp16 : unsigned(7 downto 0);
variable REG_VAR_tmp16 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_ram8_at_tmp16 := ram8_at_tmp16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_right := to_unsigned(5, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_add := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iffalse := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iftrue := to_unsigned(1, 1);
     VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_offset := resize(to_unsigned(0, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_mul := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_right := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_mul := resize(to_unsigned(1, 1), 8);
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_add := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_k := VAR_k;
     VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_left := VAR_phase;
     VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_value := ram8_at_tmp16;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue := ram8_at_tmp16;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue := ram8_at_tmp16;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse := ram8_at_tmp16;
     VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iffalse := result;
     VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_ptr := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_index := VAR_stack_index;
     VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse := t8;
     VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_address := resize(tmp16, 16);
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l748_c11_364d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l757_c11_cef8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l760_c11_169d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l742_c6_f79e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l753_c11_24df] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l745_c11_cd5f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l742_c6_f79e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l745_c11_cd5f_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l748_c11_364d_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l753_c11_24df_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l757_c11_cef8_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l760_c11_169d_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l742_c1_d064] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l760_c7_9071] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l760_c7_9071_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_cond;
     result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iftrue;
     result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output := result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l745_c7_65a3] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l742_c1_d064_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l760_c7_9071_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l745_c1_9e5b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l757_c7_5795] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond;
     result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue;
     result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output := result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l743_c12_200c] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_sp;
     set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_k;
     set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_mul;
     set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output := set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l748_c7_2112] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l745_c1_9e5b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l743_c12_200c_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l748_c1_72a3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output;

     -- t_register[uxn_opcodes_phased_h_l746_c8_d4e1] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l746_c8_d4e1_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_index;
     t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output := t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l753_c7_28d0] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond;
     result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue;
     result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output := result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l753_c7_28d0] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;
     VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l748_c1_72a3_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;
     VAR_t8_uxn_opcodes_phased_h_l746_c3_f1e4 := resize(VAR_t_register_uxn_opcodes_phased_h_l746_c8_d4e1_return_output, 16);
     VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue := VAR_t8_uxn_opcodes_phased_h_l746_c3_f1e4;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l757_c7_5795] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output;

     -- t_register[uxn_opcodes_phased_h_l749_c8_5b93] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l749_c8_5b93_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_index;
     t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output := t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l753_c1_1c15] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l748_c7_2112] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond;
     result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue;
     result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output := result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;

     -- Submodule level 5
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c7_5795_return_output;
     VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output;
     VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l753_c1_1c15_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;
     VAR_t8_uxn_opcodes_phased_h_l749_c3_4ab4 := resize(VAR_t_register_uxn_opcodes_phased_h_l749_c8_5b93_return_output, 16);
     VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue := VAR_t8_uxn_opcodes_phased_h_l749_c3_4ab4;
     -- set[uxn_opcodes_phased_h_l755_c3_0b69] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l755_c3_0b69_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l755_c3_0b69_sp <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_sp;
     set_uxn_opcodes_phased_h_l755_c3_0b69_stack_index <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_stack_index;
     set_uxn_opcodes_phased_h_l755_c3_0b69_ins <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_ins;
     set_uxn_opcodes_phased_h_l755_c3_0b69_k <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_k;
     set_uxn_opcodes_phased_h_l755_c3_0b69_mul <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_mul;
     set_uxn_opcodes_phased_h_l755_c3_0b69_add <= VAR_set_uxn_opcodes_phased_h_l755_c3_0b69_add;
     -- Outputs

     -- CAST_TO_int8_t[uxn_opcodes_phased_h_l750_c17_1f12] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_phased_h_l750_c17_1f12_return_output := CAST_TO_int8_t_uint16_t(
     VAR_t8_uxn_opcodes_phased_h_l749_c3_4ab4);

     -- result_MUX[uxn_opcodes_phased_h_l745_c7_65a3] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond;
     result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue;
     result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output := result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l748_c7_2112] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond;
     t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output := t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;

     -- peek_ram[uxn_opcodes_phased_h_l754_c19_6dee] LATENCY=0
     -- Clock enable
     peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_CLOCK_ENABLE <= VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_CLOCK_ENABLE;
     -- Inputs
     peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_address <= VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_address;
     -- Outputs
     VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output := peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l757_c1_0057] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output;

     -- Submodule level 6
     VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_right := VAR_CAST_TO_int8_t_uxn_opcodes_phased_h_l750_c17_1f12_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l757_c1_0057_return_output;
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue := VAR_peek_ram_uxn_opcodes_phased_h_l754_c19_6dee_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l745_c7_65a3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond;
     t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output := t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;

     -- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l753_c7_28d0] LATENCY=0
     -- Inputs
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_cond;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iftrue;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_iffalse;
     -- Outputs
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output := ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;

     -- put_stack[uxn_opcodes_phased_h_l758_c3_d8d5] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_sp <= VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_sp;
     put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_stack_index;
     put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_offset <= VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_offset;
     put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_value <= VAR_put_stack_uxn_opcodes_phased_h_l758_c3_d8d5_value;
     -- Outputs

     -- BIN_OP_PLUS[uxn_opcodes_phased_h_l750_c11_aeb5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_left;
     BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output := BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l742_c2_e567] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond;
     result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue;
     result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output := result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;

     -- Submodule level 7
     VAR_tmp16_uxn_opcodes_phased_h_l750_c3_ceda := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l750_c11_aeb5_return_output)),8);
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse := VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l753_c7_28d0_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;
     VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_address := resize(VAR_tmp16_uxn_opcodes_phased_h_l750_c3_ceda, 16);
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue := VAR_tmp16_uxn_opcodes_phased_h_l750_c3_ceda;
     -- peek_ram[uxn_opcodes_phased_h_l751_c19_a4da] LATENCY=0
     -- Clock enable
     peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_CLOCK_ENABLE <= VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_CLOCK_ENABLE;
     -- Inputs
     peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_address <= VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_address;
     -- Outputs
     VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output := peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output;

     -- tmp16_MUX[uxn_opcodes_phased_h_l748_c7_2112] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond;
     tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue;
     tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output := tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l742_c2_e567] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond;
     t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output := t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;

     -- Submodule level 8
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue := VAR_peek_ram_uxn_opcodes_phased_h_l751_c19_a4da_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse := VAR_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;
     -- tmp16_MUX[uxn_opcodes_phased_h_l745_c7_65a3] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond;
     tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue;
     tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output := tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;

     -- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l748_c7_2112] LATENCY=0
     -- Inputs
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_cond;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iftrue;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_iffalse;
     -- Outputs
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output := ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;

     -- Submodule level 9
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse := VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l748_c7_2112_return_output;
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse := VAR_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;
     -- tmp16_MUX[uxn_opcodes_phased_h_l742_c2_e567] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond;
     tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue;
     tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse <= VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output := tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;

     -- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l745_c7_65a3] LATENCY=0
     -- Inputs
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_cond;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iftrue;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_iffalse;
     -- Outputs
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output := ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;

     -- Submodule level 10
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse := VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l745_c7_65a3_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;
     -- ram8_at_tmp16_MUX[uxn_opcodes_phased_h_l742_c2_e567] LATENCY=0
     -- Inputs
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_cond;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iftrue;
     ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse <= VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_iffalse;
     -- Outputs
     VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output := ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;

     -- Submodule level 11
     REG_VAR_ram8_at_tmp16 := VAR_ram8_at_tmp16_MUX_uxn_opcodes_phased_h_l742_c2_e567_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_ram8_at_tmp16 <= REG_VAR_ram8_at_tmp16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     ram8_at_tmp16 <= REG_COMB_ram8_at_tmp16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
