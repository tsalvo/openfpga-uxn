-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity ora_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_64d180f1;
architecture arch of ora_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1013_c6_ac21]
signal BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal t8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal n8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1013_c2_ba69]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1026_c11_1138]
signal BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1026_c7_7735]
signal t8_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1026_c7_7735]
signal n8_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1026_c7_7735]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1026_c7_7735]
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1026_c7_7735]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1026_c7_7735]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1026_c7_7735]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1029_c11_47cd]
signal BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1029_c7_6b1a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1032_c11_01f7]
signal BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1032_c7_bb20]
signal n8_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1032_c7_bb20]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1032_c7_bb20]
signal result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1032_c7_bb20]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1032_c7_bb20]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1032_c7_bb20]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1034_c30_59a4]
signal sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1037_c21_f488]
signal BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21
BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_left,
BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_right,
BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output);

-- t8_MUX_uxn_opcodes_h_l1013_c2_ba69
t8_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- n8_MUX_uxn_opcodes_h_l1013_c2_ba69
n8_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69
result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69
result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69
result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69
result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69
result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69
result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69
result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_left,
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_right,
BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output);

-- t8_MUX_uxn_opcodes_h_l1026_c7_7735
t8_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
t8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
t8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- n8_MUX_uxn_opcodes_h_l1026_c7_7735
n8_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
n8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
n8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd
BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_left,
BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_right,
BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output);

-- t8_MUX_uxn_opcodes_h_l1029_c7_6b1a
t8_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- n8_MUX_uxn_opcodes_h_l1029_c7_6b1a
n8_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a
result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a
result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a
result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7
BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_left,
BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_right,
BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output);

-- n8_MUX_uxn_opcodes_h_l1032_c7_bb20
n8_MUX_uxn_opcodes_h_l1032_c7_bb20 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1032_c7_bb20_cond,
n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue,
n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse,
n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20
result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20
result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_cond,
result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20
result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20
result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4
sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_ins,
sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_x,
sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_y,
sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488
BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_left,
BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_right,
BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output,
 t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output,
 t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output,
 t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output,
 n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output,
 sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1018_c3_e702 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1023_c3_dd9c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1027_c3_b6b5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1036_c3_9256 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_3add_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_dcf2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_e3d6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1029_l1032_DUPLICATE_1f9e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1041_l1009_DUPLICATE_ddb0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1027_c3_b6b5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1027_c3_b6b5;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1023_c3_dd9c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1023_c3_dd9c;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1036_c3_9256 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1036_c3_9256;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1018_c3_e702 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1018_c3_e702;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_3add LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_3add_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1013_c6_ac21] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_left;
     BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output := BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_e3d6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_e3d6_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_dcf2 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_dcf2_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1034_c30_59a4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_ins;
     sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_x;
     sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output := sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1029_c11_47cd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1026_c11_1138] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_left;
     BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output := BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1029_l1032_DUPLICATE_1f9e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1029_l1032_DUPLICATE_1f9e_return_output := result.stack_address_sp_offset;

     -- BIN_OP_OR[uxn_opcodes_h_l1037_c21_f488] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_left;
     BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output := BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1032_c11_01f7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1013_c6_ac21_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1026_c11_1138_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1029_c11_47cd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1032_c11_01f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1037_c21_f488_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_dcf2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_dcf2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_dcf2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_3add_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_3add_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_3add_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_e3d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_e3d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1029_l1032_l1026_DUPLICATE_e3d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1029_l1032_DUPLICATE_1f9e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1029_l1032_DUPLICATE_1f9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1029_l1032_l1026_l1013_DUPLICATE_382d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1013_c2_ba69_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1034_c30_59a4_return_output;
     -- t8_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1032_c7_bb20] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output := result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1032_c7_bb20] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- n8_MUX[uxn_opcodes_h_l1032_c7_bb20] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1032_c7_bb20_cond <= VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_cond;
     n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue;
     n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output := n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1032_c7_bb20] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1032_c7_bb20] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1032_c7_bb20] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1032_c7_bb20_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     -- t8_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     t8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     t8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1029_c7_6b1a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1029_c7_6b1a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- t8_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- n8_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     n8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     n8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1026_c7_7735] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1026_c7_7735_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- n8_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1013_c2_ba69] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1041_l1009_DUPLICATE_ddb0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1041_l1009_DUPLICATE_ddb0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1013_c2_ba69_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1041_l1009_DUPLICATE_ddb0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1041_l1009_DUPLICATE_ddb0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
