-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity div_0CLK_622c3f98 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_622c3f98;
architecture arch of div_0CLK_622c3f98 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2023_c6_fc28]
signal BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2023_c2_213a]
signal n8_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2023_c2_213a]
signal result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2023_c2_213a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2023_c2_213a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2023_c2_213a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2023_c2_213a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2023_c2_213a]
signal t8_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2030_c11_215d]
signal BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal n8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2030_c7_fb35]
signal t8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2033_c11_2c44]
signal BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2033_c7_b2c4]
signal t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2036_c11_1a5b]
signal BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2036_c7_5f3c]
signal n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2036_c7_5f3c]
signal result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2036_c7_5f3c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2036_c7_5f3c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2036_c7_5f3c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2036_c7_5f3c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2039_c30_9415]
signal sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2042_c21_06ad]
signal BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2042_c35_cff7]
signal BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2042_c21_5234]
signal MUX_uxn_opcodes_h_l2042_c21_5234_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2042_c21_5234_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2042_c21_5234_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2042_c21_5234_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2044_c11_0939]
signal BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2044_c7_7c80]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2044_c7_7c80]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2044_c7_7c80]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28
BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_left,
BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_right,
BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output);

-- n8_MUX_uxn_opcodes_h_l2023_c2_213a
n8_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
n8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
n8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a
result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a
result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a
result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- t8_MUX_uxn_opcodes_h_l2023_c2_213a
t8_MUX_uxn_opcodes_h_l2023_c2_213a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2023_c2_213a_cond,
t8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue,
t8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse,
t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_left,
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_right,
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output);

-- n8_MUX_uxn_opcodes_h_l2030_c7_fb35
n8_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35
result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35
result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- t8_MUX_uxn_opcodes_h_l2030_c7_fb35
t8_MUX_uxn_opcodes_h_l2030_c7_fb35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond,
t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue,
t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse,
t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44
BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_left,
BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_right,
BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output);

-- n8_MUX_uxn_opcodes_h_l2033_c7_b2c4
n8_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4
result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4
result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4
result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- t8_MUX_uxn_opcodes_h_l2033_c7_b2c4
t8_MUX_uxn_opcodes_h_l2033_c7_b2c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond,
t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue,
t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse,
t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b
BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_left,
BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_right,
BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output);

-- n8_MUX_uxn_opcodes_h_l2036_c7_5f3c
n8_MUX_uxn_opcodes_h_l2036_c7_5f3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond,
n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue,
n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse,
n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c
result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c
result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c
result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2039_c30_9415
sp_relative_shift_uxn_opcodes_h_l2039_c30_9415 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_ins,
sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_x,
sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_y,
sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad
BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_left,
BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_right,
BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7
BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_left,
BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_right,
BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output);

-- MUX_uxn_opcodes_h_l2042_c21_5234
MUX_uxn_opcodes_h_l2042_c21_5234 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2042_c21_5234_cond,
MUX_uxn_opcodes_h_l2042_c21_5234_iftrue,
MUX_uxn_opcodes_h_l2042_c21_5234_iffalse,
MUX_uxn_opcodes_h_l2042_c21_5234_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939
BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_left,
BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_right,
BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80
result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80
result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80
result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output,
 n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output,
 n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output,
 n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output,
 n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output,
 MUX_uxn_opcodes_h_l2042_c21_5234_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2027_c3_8782 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2031_c3_4672 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2041_c3_23b1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2042_c21_5234_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2042_c21_5234_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2042_c21_5234_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2042_c21_5234_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2045_c3_90ff : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2036_l2033_DUPLICATE_a871_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2050_l2019_DUPLICATE_fc3b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2031_c3_4672 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2031_c3_4672;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2042_c21_5234_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2027_c3_8782 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2027_c3_8782;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2045_c3_90ff := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2045_c3_90ff;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2041_c3_23b1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2041_c3_23b1;
     VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2023_c6_fc28] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_left;
     BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output := BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2030_c11_215d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2044_c11_0939] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_left;
     BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output := BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2033_c11_2c44] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_left;
     BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output := BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2042_c21_06ad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_left;
     BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output := BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2036_c11_1a5b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19_return_output := result.is_opc_done;

     -- BIN_OP_DIV[uxn_opcodes_h_l2042_c35_cff7] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_left;
     BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output := BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2039_c30_9415] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_ins;
     sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_x;
     sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output := sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2036_l2033_DUPLICATE_a871 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2036_l2033_DUPLICATE_a871_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2042_c21_5234_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2042_c35_cff7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2023_c6_fc28_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_215d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2033_c11_2c44_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2036_c11_1a5b_return_output;
     VAR_MUX_uxn_opcodes_h_l2042_c21_5234_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2042_c21_06ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2044_c11_0939_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_d024_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2036_l2030_l2044_l2033_DUPLICATE_2b19_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2030_l2044_l2033_l2023_DUPLICATE_7e05_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2036_l2033_DUPLICATE_a871_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2036_l2033_DUPLICATE_a871_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2036_l2030_l2033_l2023_DUPLICATE_a111_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2039_c30_9415_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2044_c7_7c80] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2044_c7_7c80] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2036_c7_5f3c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2036_c7_5f3c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond;
     n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue;
     n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output := n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2044_c7_7c80] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output;

     -- MUX[uxn_opcodes_h_l2042_c21_5234] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2042_c21_5234_cond <= VAR_MUX_uxn_opcodes_h_l2042_c21_5234_cond;
     MUX_uxn_opcodes_h_l2042_c21_5234_iftrue <= VAR_MUX_uxn_opcodes_h_l2042_c21_5234_iftrue;
     MUX_uxn_opcodes_h_l2042_c21_5234_iffalse <= VAR_MUX_uxn_opcodes_h_l2042_c21_5234_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2042_c21_5234_return_output := MUX_uxn_opcodes_h_l2042_c21_5234_return_output;

     -- t8_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue := VAR_MUX_uxn_opcodes_h_l2042_c21_5234_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2044_c7_7c80_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- n8_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- t8_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2036_c7_5f3c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2036_c7_5f3c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2036_c7_5f3c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2036_c7_5f3c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2036_c7_5f3c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- n8_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- t8_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     t8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     t8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2033_c7_b2c4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output := result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2033_c7_b2c4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- n8_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     n8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     n8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2030_c7_fb35] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2030_c7_fb35_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2023_c2_213a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2050_l2019_DUPLICATE_fc3b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2050_l2019_DUPLICATE_fc3b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2023_c2_213a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2023_c2_213a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2050_l2019_DUPLICATE_fc3b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2050_l2019_DUPLICATE_fc3b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
