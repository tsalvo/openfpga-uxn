-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_367c]
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2639_c2_969a]
signal n8_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_969a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2639_c2_969a]
signal l8_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2639_c2_969a]
signal t8_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_6f6e]
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2652_c7_4208]
signal n8_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_4208]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_4208]
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_4208]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_4208]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_4208]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2652_c7_4208]
signal l8_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2652_c7_4208]
signal t8_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_eae3]
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal n8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal l8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2655_c7_ca00]
signal t8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_555e]
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2659_c7_1424]
signal n8_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_1424]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_1424]
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_1424]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_1424]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_1424]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2659_c7_1424]
signal l8_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2661_c30_4e35]
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_8714]
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_12e7]
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_12e7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_12e7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_12e7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2666_c7_12e7]
signal l8_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_e0ed]
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_2bcf]
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_2bcf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_2bcf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_left,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_right,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output);

-- n8_MUX_uxn_opcodes_h_l2639_c2_969a
n8_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
n8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
n8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- l8_MUX_uxn_opcodes_h_l2639_c2_969a
l8_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
l8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
l8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- t8_MUX_uxn_opcodes_h_l2639_c2_969a
t8_MUX_uxn_opcodes_h_l2639_c2_969a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2639_c2_969a_cond,
t8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue,
t8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse,
t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_left,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_right,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output);

-- n8_MUX_uxn_opcodes_h_l2652_c7_4208
n8_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
n8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
n8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- l8_MUX_uxn_opcodes_h_l2652_c7_4208
l8_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
l8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
l8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- t8_MUX_uxn_opcodes_h_l2652_c7_4208
t8_MUX_uxn_opcodes_h_l2652_c7_4208 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2652_c7_4208_cond,
t8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue,
t8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse,
t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_left,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_right,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output);

-- n8_MUX_uxn_opcodes_h_l2655_c7_ca00
n8_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- l8_MUX_uxn_opcodes_h_l2655_c7_ca00
l8_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- t8_MUX_uxn_opcodes_h_l2655_c7_ca00
t8_MUX_uxn_opcodes_h_l2655_c7_ca00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond,
t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue,
t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse,
t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_left,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_right,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output);

-- n8_MUX_uxn_opcodes_h_l2659_c7_1424
n8_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
n8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
n8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- l8_MUX_uxn_opcodes_h_l2659_c7_1424
l8_MUX_uxn_opcodes_h_l2659_c7_1424 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2659_c7_1424_cond,
l8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue,
l8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse,
l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35
sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_ins,
sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_x,
sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_y,
sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_left,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_right,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output);

-- l8_MUX_uxn_opcodes_h_l2666_c7_12e7
l8_MUX_uxn_opcodes_h_l2666_c7_12e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2666_c7_12e7_cond,
l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue,
l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse,
l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_left,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_right,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output,
 n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output,
 n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output,
 n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output,
 n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output,
 sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output,
 l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_5827 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_01f3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_c530 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_ed0b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_1d7f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_9d28 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_a4d5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_8fb0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_2bcf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_2dae_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_7ecb_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2678_l2635_DUPLICATE_8492_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_5827 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_5827;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_a4d5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_a4d5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_c530 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_c530;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_01f3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_01f3;
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_8fb0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_8fb0;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_ed0b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_ed0b;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_9d28 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_9d28;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_1d7f := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_1d7f;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_367c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2672_c7_2bcf] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_2bcf_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2661_c30_4e35] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_ins;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_x;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output := sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_969a_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_6f6e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_eae3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_969a_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_555e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_969a_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_2dae LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_2dae_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_e0ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_7ecb LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_7ecb_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_8714] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_left;
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output := BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_969a_return_output := result.is_ram_write;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_367c_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_6f6e_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_eae3_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_555e_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_8714_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_e0ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_7ecb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_7ecb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_7ecb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_3a52_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_2dae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_2dae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_2dae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_1e3a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_969a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_969a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_969a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_969a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_2bcf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_4e35_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_12e7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_2bcf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output;

     -- l8_MUX[uxn_opcodes_h_l2666_c7_12e7] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2666_c7_12e7_cond <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_cond;
     l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue;
     l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output := l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_2bcf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_2bcf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output;

     -- t8_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     n8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     n8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_2bcf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_12e7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_12e7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- t8_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     t8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     t8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_12e7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;

     -- l8_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     l8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     l8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_12e7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- l8_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- n8_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     n8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     n8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_1424] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output := result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;

     -- t8_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     t8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     t8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_1424_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;
     -- l8_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     l8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     l8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_ca00] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- n8_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     n8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     n8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_ca00_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_4208] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;

     -- l8_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     l8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     l8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_4208_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_969a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2678_l2635_DUPLICATE_8492 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2678_l2635_DUPLICATE_8492_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_969a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_969a_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2678_l2635_DUPLICATE_8492_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2678_l2635_DUPLICATE_8492_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
