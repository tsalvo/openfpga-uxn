-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity div_0CLK_4e24eea7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_4e24eea7;
architecture arch of div_0CLK_4e24eea7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2056_c6_2e29]
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal n8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal t8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c2_9c06]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_318e]
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal n8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal t8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_dad5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2072_c11_3fcd]
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal n8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal t8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2072_c7_92a0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2075_c11_2fdd]
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2075_c7_887b]
signal n8_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2075_c7_887b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2075_c7_887b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2075_c7_887b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2075_c7_887b]
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2075_c7_887b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2077_c30_d450]
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2080_c21_d9ee]
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2080_c35_fd14]
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2080_c21_ac7f]
signal MUX_uxn_opcodes_h_l2080_c21_ac7f_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_ac7f_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_ac7f_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_left,
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_right,
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output);

-- n8_MUX_uxn_opcodes_h_l2056_c2_9c06
n8_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- t8_MUX_uxn_opcodes_h_l2056_c2_9c06
t8_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_left,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_right,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output);

-- n8_MUX_uxn_opcodes_h_l2069_c7_dad5
n8_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- t8_MUX_uxn_opcodes_h_l2069_c7_dad5
t8_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_left,
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_right,
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output);

-- n8_MUX_uxn_opcodes_h_l2072_c7_92a0
n8_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- t8_MUX_uxn_opcodes_h_l2072_c7_92a0
t8_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_left,
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_right,
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output);

-- n8_MUX_uxn_opcodes_h_l2075_c7_887b
n8_MUX_uxn_opcodes_h_l2075_c7_887b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2075_c7_887b_cond,
n8_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue,
n8_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse,
n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2077_c30_d450
sp_relative_shift_uxn_opcodes_h_l2077_c30_d450 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_ins,
sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_x,
sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_y,
sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_left,
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_right,
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_371b3c10 port map (
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_left,
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_right,
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output);

-- MUX_uxn_opcodes_h_l2080_c21_ac7f
MUX_uxn_opcodes_h_l2080_c21_ac7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2080_c21_ac7f_cond,
MUX_uxn_opcodes_h_l2080_c21_ac7f_iftrue,
MUX_uxn_opcodes_h_l2080_c21_ac7f_iffalse,
MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output,
 n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output,
 n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output,
 n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output,
 n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output,
 MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_4a98 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_dafd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_1623 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_4a82 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_513d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_b3ab_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_daac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_b66f_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2084_l2052_DUPLICATE_4801_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_4a98 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_4a98;
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_dafd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_dafd;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_4a82 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_4a82;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_1623 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_1623;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_b66f LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_b66f_return_output := result.stack_address_sp_offset;

     -- BIN_OP_DIV[uxn_opcodes_h_l2080_c35_fd14] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_left;
     BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output := BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_b3ab LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_b3ab_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2072_c11_3fcd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2056_c6_2e29] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_left;
     BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output := BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2075_c11_2fdd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2077_c30_d450] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_ins;
     sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_x;
     sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output := sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_318e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_daac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_daac_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_513d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_513d_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2080_c21_d9ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_fd14_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_2e29_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_318e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_3fcd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_2fdd_return_output;
     VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_d9ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_513d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_513d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_513d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_b3ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_b3ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_b3ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_daac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_daac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2069_l2075_DUPLICATE_daac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_b66f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_b66f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2056_l2072_l2069_l2075_DUPLICATE_92f7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_9c06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_d450_return_output;
     -- t8_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2075_c7_887b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2075_c7_887b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;

     -- MUX[uxn_opcodes_h_l2080_c21_ac7f] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2080_c21_ac7f_cond <= VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_cond;
     MUX_uxn_opcodes_h_l2080_c21_ac7f_iftrue <= VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_iftrue;
     MUX_uxn_opcodes_h_l2080_c21_ac7f_iffalse <= VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output := MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2075_c7_887b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;

     -- n8_MUX[uxn_opcodes_h_l2075_c7_887b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2075_c7_887b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_cond;
     n8_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue;
     n8_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output := n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2075_c7_887b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue := VAR_MUX_uxn_opcodes_h_l2080_c21_ac7f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2075_c7_887b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- n8_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_887b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2072_c7_92a0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;

     -- n8_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- t8_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_92a0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_dad5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- n8_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_dad5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2056_c2_9c06] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output := result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2084_l2052_DUPLICATE_4801 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2084_l2052_DUPLICATE_4801_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_9c06_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2084_l2052_DUPLICATE_4801_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2084_l2052_DUPLICATE_4801_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
