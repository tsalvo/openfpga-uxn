-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_64d180f1;
architecture arch of eor_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1093_c6_e06a]
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal n8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1093_c2_7b97]
signal t8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1106_c11_abb8]
signal BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal n8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1106_c7_bda4]
signal t8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1109_c11_ab88]
signal BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal n8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1109_c7_4f87]
signal t8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1112_c11_3285]
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1112_c7_8d6d]
signal n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1112_c7_8d6d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1112_c7_8d6d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1112_c7_8d6d]
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1112_c7_8d6d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1112_c7_8d6d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1114_c30_2c1f]
signal sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1117_c21_4046]
signal BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_left,
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_right,
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output);

-- n8_MUX_uxn_opcodes_h_l1093_c2_7b97
n8_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97
result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97
result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97
result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- t8_MUX_uxn_opcodes_h_l1093_c2_7b97
t8_MUX_uxn_opcodes_h_l1093_c2_7b97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond,
t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue,
t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse,
t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8
BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_left,
BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_right,
BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output);

-- n8_MUX_uxn_opcodes_h_l1106_c7_bda4
n8_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4
result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4
result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4
result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- t8_MUX_uxn_opcodes_h_l1106_c7_bda4
t8_MUX_uxn_opcodes_h_l1106_c7_bda4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond,
t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue,
t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse,
t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88
BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_left,
BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_right,
BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output);

-- n8_MUX_uxn_opcodes_h_l1109_c7_4f87
n8_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87
result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87
result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87
result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87
result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- t8_MUX_uxn_opcodes_h_l1109_c7_4f87
t8_MUX_uxn_opcodes_h_l1109_c7_4f87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond,
t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue,
t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse,
t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_left,
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_right,
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output);

-- n8_MUX_uxn_opcodes_h_l1112_c7_8d6d
n8_MUX_uxn_opcodes_h_l1112_c7_8d6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond,
n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue,
n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse,
n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f
sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_ins,
sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_x,
sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_y,
sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046
BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046 : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_left,
BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_right,
BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output,
 n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output,
 n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output,
 n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output,
 n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output,
 sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1098_c3_2994 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1103_c3_22f7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1107_c3_7176 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_95b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_f078_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1d5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1c0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1112_l1109_DUPLICATE_1525_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1089_l1121_DUPLICATE_87f1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_95b0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_95b0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1103_c3_22f7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1103_c3_22f7;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1107_c3_7176 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1107_c3_7176;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1098_c3_2994 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1098_c3_2994;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1112_l1109_DUPLICATE_1525 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1112_l1109_DUPLICATE_1525_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1d5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1d5_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1106_c11_abb8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1109_c11_ab88] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_left;
     BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output := BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1c0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1c0_return_output := result.is_stack_write;

     -- BIN_OP_XOR[uxn_opcodes_h_l1117_c21_4046] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_left;
     BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output := BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1114_c30_2c1f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_ins;
     sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_x;
     sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output := sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1093_c6_e06a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1112_c11_3285] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_left;
     BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output := BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_f078 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_f078_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_e06a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1106_c11_abb8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1109_c11_ab88_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_3285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1117_c21_4046_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_f078_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_f078_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1106_l1109_l1112_DUPLICATE_a1c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1112_l1109_DUPLICATE_1525_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1112_l1109_DUPLICATE_1525_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1106_l1109_l1112_l1093_DUPLICATE_d645_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1093_c2_7b97_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1114_c30_2c1f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1112_c7_8d6d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1112_c7_8d6d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1112_c7_8d6d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;

     -- n8_MUX[uxn_opcodes_h_l1112_c7_8d6d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond;
     n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue;
     n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output := n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1112_c7_8d6d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1112_c7_8d6d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- t8_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_8d6d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- n8_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- t8_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1109_c7_4f87] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1109_c7_4f87_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     -- n8_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1106_c7_bda4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1106_c7_bda4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- n8_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c2_7b97] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1089_l1121_DUPLICATE_87f1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1089_l1121_DUPLICATE_87f1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1093_c2_7b97_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1089_l1121_DUPLICATE_87f1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1089_l1121_DUPLICATE_87f1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
