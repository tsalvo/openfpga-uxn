-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity rot_0CLK_57104a4d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_57104a4d;
architecture arch of rot_0CLK_57104a4d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2602_c6_973a]
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal n8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal l8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2602_c2_f22e]
signal t8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2609_c11_fcb1]
signal BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2609_c7_9698]
signal n8_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2609_c7_9698]
signal l8_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2609_c7_9698]
signal result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2609_c7_9698]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2609_c7_9698]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2609_c7_9698]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2609_c7_9698]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2609_c7_9698]
signal t8_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2612_c11_c403]
signal BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal n8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal l8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2612_c7_d89e]
signal t8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2616_c11_56ca]
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2616_c7_2c9c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2619_c30_5988]
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_5414]
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2624_c7_21b9]
signal l8_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2624_c7_21b9]
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_21b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_21b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2624_c7_21b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2624_c7_21b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2630_c11_befe]
signal BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2630_c7_cede]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2630_c7_cede]
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2630_c7_cede]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2630_c7_cede]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2634_c11_3754]
signal BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2634_c7_8f85]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2634_c7_8f85]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_left,
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_right,
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output);

-- n8_MUX_uxn_opcodes_h_l2602_c2_f22e
n8_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- l8_MUX_uxn_opcodes_h_l2602_c2_f22e
l8_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- t8_MUX_uxn_opcodes_h_l2602_c2_f22e
t8_MUX_uxn_opcodes_h_l2602_c2_f22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond,
t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue,
t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse,
t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_left,
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_right,
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output);

-- n8_MUX_uxn_opcodes_h_l2609_c7_9698
n8_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
n8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
n8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- l8_MUX_uxn_opcodes_h_l2609_c7_9698
l8_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
l8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
l8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698
result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- t8_MUX_uxn_opcodes_h_l2609_c7_9698
t8_MUX_uxn_opcodes_h_l2609_c7_9698 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2609_c7_9698_cond,
t8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue,
t8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse,
t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403
BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_left,
BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_right,
BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output);

-- n8_MUX_uxn_opcodes_h_l2612_c7_d89e
n8_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- l8_MUX_uxn_opcodes_h_l2612_c7_d89e
l8_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e
result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e
result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e
result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- t8_MUX_uxn_opcodes_h_l2612_c7_d89e
t8_MUX_uxn_opcodes_h_l2612_c7_d89e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond,
t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue,
t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse,
t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_left,
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_right,
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output);

-- n8_MUX_uxn_opcodes_h_l2616_c7_2c9c
n8_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- l8_MUX_uxn_opcodes_h_l2616_c7_2c9c
l8_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2619_c30_5988
sp_relative_shift_uxn_opcodes_h_l2619_c30_5988 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_ins,
sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_x,
sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_y,
sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_left,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_right,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output);

-- l8_MUX_uxn_opcodes_h_l2624_c7_21b9
l8_MUX_uxn_opcodes_h_l2624_c7_21b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2624_c7_21b9_cond,
l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue,
l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse,
l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_left,
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_right,
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_cond,
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_left,
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_right,
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output,
 n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output,
 n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output,
 n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output,
 n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output,
 l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2606_c3_5825 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2610_c3_2a46 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2613_c3_dc79 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_60b5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2627_c3_dfc4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2626_c3_70c4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2631_c3_7e07 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2630_c7_cede_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2598_l2639_DUPLICATE_32da_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2631_c3_7e07 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2631_c3_7e07;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_60b5 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_60b5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_right := to_unsigned(6, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2610_c3_2a46 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2610_c3_2a46;
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2613_c3_dc79 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2613_c3_dc79;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2626_c3_70c4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2626_c3_70c4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2627_c3_dfc4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2627_c3_dfc4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2606_c3_5825 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2606_c3_5825;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l2619_c30_5988] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_ins;
     sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_x;
     sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output := sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2630_c7_cede] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2630_c7_cede_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2612_c11_c403] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_left;
     BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output := BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2634_c11_3754] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_left;
     BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output := BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2630_c11_befe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_left;
     BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output := BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2609_c11_fcb1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_5414] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_left;
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output := BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2616_c11_56ca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_left;
     BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output := BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2602_c6_973a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_973a_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_fcb1_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2612_c11_c403_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_56ca_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_5414_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_befe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_3754_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2609_l2624_l2612_l2602_DUPLICATE_fec1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2634_l2630_l2624_l2616_l2612_DUPLICATE_0be5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2602_l2634_l2630_l2624_l2612_DUPLICATE_6bee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2609_l2612_l2630_l2602_DUPLICATE_9744_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2630_c7_cede_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_5988_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2624_c7_21b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2634_c7_8f85] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2634_c7_8f85] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output;

     -- t8_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2630_c7_cede] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;

     -- n8_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2630_c7_cede] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output := result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;

     -- l8_MUX[uxn_opcodes_h_l2624_c7_21b9] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2624_c7_21b9_cond <= VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_cond;
     l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue;
     l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output := l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_8f85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2630_c7_cede] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2630_c7_cede] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;

     -- l8_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2624_c7_21b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     t8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     t8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2624_c7_21b9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_cede_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_21b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- l8_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     n8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     n8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_21b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_21b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;
     -- n8_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- l8_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     l8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     l8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2616_c7_2c9c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_2c9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- l8_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2612_c7_d89e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2612_c7_d89e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2609_c7_9698] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_9698_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2602_c2_f22e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2598_l2639_DUPLICATE_32da LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2598_l2639_DUPLICATE_32da_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_f22e_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2598_l2639_DUPLICATE_32da_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2598_l2639_DUPLICATE_32da_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
