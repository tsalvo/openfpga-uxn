-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sth_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_85d5529e;
architecture arch of sth_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2542_c6_1994]
signal BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2542_c1_d04e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2542_c2_40e2]
signal t8_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2543_c3_7f25[uxn_opcodes_h_l2543_c3_7f25]
signal printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2547_c11_1b38]
signal BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2547_c7_8716]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2547_c7_8716]
signal t8_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2550_c11_90bb]
signal BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2550_c7_f7e3]
signal t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2553_c30_4c37]
signal sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2555_c11_e3f3]
signal BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2555_c7_4278]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2562_c11_864e]
signal BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2562_c7_5cd2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2562_c7_5cd2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2562_c7_5cd2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2562_c7_5cd2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_78f9( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994
BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_left,
BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_right,
BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2
result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2
result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2
result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2
result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- t8_MUX_uxn_opcodes_h_l2542_c2_40e2
t8_MUX_uxn_opcodes_h_l2542_c2_40e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2542_c2_40e2_cond,
t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue,
t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse,
t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

-- printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25
printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25 : entity work.printf_uxn_opcodes_h_l2543_c3_7f25_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38
BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_left,
BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_right,
BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716
result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716
result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716
result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716
result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716
result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- t8_MUX_uxn_opcodes_h_l2547_c7_8716
t8_MUX_uxn_opcodes_h_l2547_c7_8716 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2547_c7_8716_cond,
t8_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue,
t8_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse,
t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb
BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_left,
BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_right,
BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- t8_MUX_uxn_opcodes_h_l2550_c7_f7e3
t8_MUX_uxn_opcodes_h_l2550_c7_f7e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond,
t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue,
t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse,
t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37
sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_ins,
sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_x,
sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_y,
sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3
BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_left,
BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_right,
BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278
result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278
result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278
result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278
result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278
result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e
BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_left,
BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_right,
BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2
result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2
result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2
result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output,
 sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2544_c3_9e60 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2548_c3_9e53 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2559_c3_2f37 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2557_c3_8e51 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_DUPLICATE_4195_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2550_l2555_DUPLICATE_493a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_78f9_uxn_opcodes_h_l2569_l2538_DUPLICATE_82f1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2544_c3_9e60 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2544_c3_9e60;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2559_c3_2f37 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2559_c3_2f37;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2557_c3_8e51 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2557_c3_8e51;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2548_c3_9e53 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2548_c3_9e53;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2562_c11_864e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2553_c30_4c37] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_ins;
     sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_x;
     sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output := sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2555_c11_e3f3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2550_c11_90bb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2542_c6_1994] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_left;
     BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output := BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_DUPLICATE_4195 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_DUPLICATE_4195_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2547_c11_1b38] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_left;
     BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output := BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2550_l2555_DUPLICATE_493a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2550_l2555_DUPLICATE_493a_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2542_c6_1994_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2547_c11_1b38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2550_c11_90bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2555_c11_e3f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2562_c11_864e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_DUPLICATE_4195_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_DUPLICATE_4195_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_DUPLICATE_4195_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2550_l2555_l2547_l2562_DUPLICATE_90d5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2542_l2555_l2547_l2562_DUPLICATE_5e24_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_88d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2550_l2542_l2547_l2562_DUPLICATE_ee58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2550_l2555_DUPLICATE_493a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2550_l2555_DUPLICATE_493a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2550_l2542_l2555_l2547_DUPLICATE_4b35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2553_c30_4c37_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2562_c7_5cd2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2562_c7_5cd2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2542_c1_d04e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2562_c7_5cd2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2562_c7_5cd2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2542_c1_d04e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2562_c7_5cd2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     -- printf_uxn_opcodes_h_l2543_c3_7f25[uxn_opcodes_h_l2543_c3_7f25] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2543_c3_7f25_uxn_opcodes_h_l2543_c3_7f25_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- t8_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     t8_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     t8_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2555_c7_4278] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2555_c7_4278_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- t8_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2550_c7_f7e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2550_c7_f7e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2547_c7_8716] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2547_c7_8716_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2542_c2_40e2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_78f9_uxn_opcodes_h_l2569_l2538_DUPLICATE_82f1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_78f9_uxn_opcodes_h_l2569_l2538_DUPLICATE_82f1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_78f9(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2542_c2_40e2_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_78f9_uxn_opcodes_h_l2569_l2538_DUPLICATE_82f1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_78f9_uxn_opcodes_h_l2569_l2538_DUPLICATE_82f1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
