-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity str1_0CLK_1e72bf9c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end str1_0CLK_1e72bf9c;
architecture arch of str1_0CLK_1e72bf9c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1687_c6_d3d2]
signal BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal n8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1687_c2_10fe]
signal t8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1700_c11_a611]
signal BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal n8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1700_c7_da8f]
signal t8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1703_c11_041a]
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1703_c7_7f2b]
signal t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1706_c11_6d9e]
signal BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1706_c7_c0bc]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1706_c7_c0bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1706_c7_c0bc]
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1706_c7_c0bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1706_c7_c0bc]
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l1706_c7_c0bc]
signal n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1708_c30_523c]
signal sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output : signed(3 downto 0);

-- u16_add_u8_as_i8[uxn_opcodes_h_l1710_c22_beab]
signal u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u16 : unsigned(15 downto 0);
signal u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u8 : unsigned(7 downto 0);
signal u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output : unsigned(15 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_ram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.u16_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2
BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_left,
BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_right,
BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe
result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe
result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe
result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe
result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe
result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe
result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe
result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe
result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- n8_MUX_uxn_opcodes_h_l1687_c2_10fe
n8_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- t8_MUX_uxn_opcodes_h_l1687_c2_10fe
t8_MUX_uxn_opcodes_h_l1687_c2_10fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond,
t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue,
t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse,
t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_left,
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_right,
BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f
result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- n8_MUX_uxn_opcodes_h_l1700_c7_da8f
n8_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- t8_MUX_uxn_opcodes_h_l1700_c7_da8f
t8_MUX_uxn_opcodes_h_l1700_c7_da8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond,
t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue,
t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse,
t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_left,
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_right,
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b
result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- n8_MUX_uxn_opcodes_h_l1703_c7_7f2b
n8_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- t8_MUX_uxn_opcodes_h_l1703_c7_7f2b
t8_MUX_uxn_opcodes_h_l1703_c7_7f2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond,
t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue,
t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse,
t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_left,
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_right,
BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc
result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond,
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output);

-- n8_MUX_uxn_opcodes_h_l1706_c7_c0bc
n8_MUX_uxn_opcodes_h_l1706_c7_c0bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond,
n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue,
n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse,
n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1708_c30_523c
sp_relative_shift_uxn_opcodes_h_l1708_c30_523c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_ins,
sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_x,
sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_y,
sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output);

-- u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab
u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab : entity work.u16_add_u8_as_i8_0CLK_e595f783 port map (
u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u16,
u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u8,
u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output,
 n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output,
 sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output,
 u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1697_c3_3186 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1692_c3_daa4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1701_c3_0d9b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1700_c7_da8f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output : signed(3 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u16 : unsigned(15 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u8 : unsigned(7 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_ecb1_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f6c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f82_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1683_l1715_DUPLICATE_7535_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1697_c3_3186 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1697_c3_3186;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1692_c3_daa4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1692_c3_daa4;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1701_c3_0d9b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1701_c3_0d9b;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse := n8;
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u16 := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := t8;
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u8 := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_ecb1 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_ecb1_return_output := result.sp_relative_shift;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1687_c6_d3d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc_return_output := result.u8_value;

     -- u16_add_u8_as_i8[uxn_opcodes_h_l1710_c22_beab] LATENCY=0
     -- Inputs
     u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u16 <= VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u16;
     u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u8 <= VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_u8;
     -- Outputs
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output := u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1700_c11_a611] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_left;
     BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output := BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f82 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f82_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f6c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f6c_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1706_c11_6d9e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1708_c30_523c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_ins;
     sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_x;
     sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output := sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1703_c11_041a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1700_c7_da8f_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1687_c6_d3d2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1700_c11_a611_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_041a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1706_c11_6d9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_ecb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_ecb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_ecb1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_ccf0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f6c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f82_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f82_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1703_l1706_l1700_DUPLICATE_5f82_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1703_l1687_l1706_l1700_DUPLICATE_66dc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1687_c2_10fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1708_c30_523c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue := VAR_u16_add_u8_as_i8_uxn_opcodes_h_l1710_c22_beab_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1706_c7_c0bc] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1706_c7_c0bc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output := result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;

     -- t8_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- n8_MUX[uxn_opcodes_h_l1706_c7_c0bc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond <= VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond;
     n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue;
     n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output := n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1706_c7_c0bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1706_c7_c0bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1706_c7_c0bc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1706_c7_c0bc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     -- t8_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- n8_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1703_c7_7f2b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_7f2b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     -- n8_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1700_c7_da8f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1700_c7_da8f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- n8_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1687_c2_10fe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1683_l1715_DUPLICATE_7535 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1683_l1715_DUPLICATE_7535_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1687_c2_10fe_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1683_l1715_DUPLICATE_7535_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l1683_l1715_DUPLICATE_7535_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
