-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity dup2_0CLK_0d289325 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end dup2_0CLK_0d289325;
architecture arch of dup2_0CLK_0d289325 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2483_c6_372b]
signal BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2483_c2_3b43]
signal t16_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2491_c11_7b0f]
signal BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2491_c7_dad5]
signal t16_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2493_c30_771e]
signal sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2495_c11_c991]
signal BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2495_c7_4b7d]
signal t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2502_c11_3ab5]
signal BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2502_c7_c1d9]
signal result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2502_c7_c1d9]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2502_c7_c1d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2502_c7_c1d9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2502_c7_c1d9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2506_c11_83fb]
signal BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2506_c7_7cf7]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2506_c7_7cf7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2506_c7_7cf7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b
BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_left,
BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_right,
BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43
result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43
result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43
result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43
result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43
result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- t16_MUX_uxn_opcodes_h_l2483_c2_3b43
t16_MUX_uxn_opcodes_h_l2483_c2_3b43 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2483_c2_3b43_cond,
t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue,
t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse,
t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_left,
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_right,
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5
result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5
result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- t16_MUX_uxn_opcodes_h_l2491_c7_dad5
t16_MUX_uxn_opcodes_h_l2491_c7_dad5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2491_c7_dad5_cond,
t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue,
t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse,
t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2493_c30_771e
sp_relative_shift_uxn_opcodes_h_l2493_c30_771e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_ins,
sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_x,
sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_y,
sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_left,
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_right,
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d
result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d
result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- t16_MUX_uxn_opcodes_h_l2495_c7_4b7d
t16_MUX_uxn_opcodes_h_l2495_c7_4b7d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond,
t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue,
t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse,
t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5
BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_left,
BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_right,
BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9
result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond,
result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9
result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9
result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb
BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_left,
BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_right,
BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7
result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7
result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output,
 sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2488_c3_23a9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2499_c3_ab7e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2503_c3_846b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2495_l2483_DUPLICATE_6c65_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2483_l2502_l2491_DUPLICATE_b830_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2483_l2491_DUPLICATE_69dd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2502_l2491_DUPLICATE_d6df_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2512_l2479_DUPLICATE_0122_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2499_c3_ab7e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2499_c3_ab7e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2488_c3_23a9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2488_c3_23a9;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2503_c3_846b := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2503_c3_846b;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_left := VAR_phase;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2495_c11_c991] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_left;
     BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output := BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2502_c11_3ab5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2502_l2491_DUPLICATE_d6df LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2502_l2491_DUPLICATE_d6df_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2483_l2491_DUPLICATE_69dd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2483_l2491_DUPLICATE_69dd_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2506_c11_83fb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2483_l2502_l2491_DUPLICATE_b830 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2483_l2502_l2491_DUPLICATE_b830_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2495_l2483_DUPLICATE_6c65 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2495_l2483_DUPLICATE_6c65_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2483_c6_372b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2493_c30_771e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_ins;
     sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_x;
     sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output := sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2491_c11_7b0f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2483_c6_372b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_7b0f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_c991_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2502_c11_3ab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2506_c11_83fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2483_l2491_DUPLICATE_69dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2483_l2491_DUPLICATE_69dd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2483_l2502_l2491_DUPLICATE_b830_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2483_l2502_l2491_DUPLICATE_b830_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2483_l2502_l2491_DUPLICATE_b830_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_4c9c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2495_l2483_DUPLICATE_6c65_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2495_l2483_DUPLICATE_6c65_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2495_l2502_l2491_l2506_DUPLICATE_f2f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2483_l2502_l2491_l2506_DUPLICATE_b4b7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2502_l2491_DUPLICATE_d6df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2502_l2491_DUPLICATE_d6df_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2493_c30_771e_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2506_c7_7cf7] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2502_c7_c1d9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2502_c7_c1d9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output := result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2506_c7_7cf7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output;

     -- t16_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2506_c7_7cf7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2506_c7_7cf7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2502_c7_c1d9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2502_c7_c1d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;

     -- t16_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2502_c7_c1d9] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2502_c7_c1d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- t16_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2495_c7_4b7d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_4b7d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2491_c7_dad5] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_dad5_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2483_c2_3b43] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2512_l2479_DUPLICATE_0122 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2512_l2479_DUPLICATE_0122_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2483_c2_3b43_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2512_l2479_DUPLICATE_0122_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2512_l2479_DUPLICATE_0122_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
