-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ldz_0CLK_46731a7b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_46731a7b;
architecture arch of ldz_0CLK_46731a7b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1523_c6_295a]
signal BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1523_c1_0ab8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1523_c2_f166]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1523_c2_f166]
signal tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1523_c2_f166]
signal t8_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1524_c3_43be[uxn_opcodes_h_l1524_c3_43be]
signal printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1528_c11_7086]
signal BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1528_c7_9392]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1528_c7_9392]
signal tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1528_c7_9392]
signal t8_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1531_c11_f311]
signal BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1531_c7_5c81]
signal t8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1534_c30_60ef]
signal sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1537_c11_8e86]
signal BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1537_c7_b42c]
signal tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1541_c11_d466]
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1541_c7_94b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1541_c7_94b3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1541_c7_94b3]
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1541_c7_94b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1541_c7_94b3]
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1547_c11_8f7e]
signal BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1547_c7_cd18]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1547_c7_cd18]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_284d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u16_value := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a
BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_left,
BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_right,
BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166
result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166
result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1523_c2_f166
tmp8_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- t8_MUX_uxn_opcodes_h_l1523_c2_f166
t8_MUX_uxn_opcodes_h_l1523_c2_f166 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1523_c2_f166_cond,
t8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue,
t8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse,
t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

-- printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be
printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be : entity work.printf_uxn_opcodes_h_l1524_c3_43be_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086
BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_left,
BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_right,
BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392
result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392
result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392
result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392
result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392
result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392
result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1528_c7_9392
tmp8_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- t8_MUX_uxn_opcodes_h_l1528_c7_9392
t8_MUX_uxn_opcodes_h_l1528_c7_9392 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1528_c7_9392_cond,
t8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue,
t8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse,
t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311
BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_left,
BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_right,
BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81
result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81
result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81
result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81
result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81
result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81
result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81
tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- t8_MUX_uxn_opcodes_h_l1531_c7_5c81
t8_MUX_uxn_opcodes_h_l1531_c7_5c81 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond,
t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue,
t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse,
t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef
sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_ins,
sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_x,
sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_y,
sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86
BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_left,
BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_right,
BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c
result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c
result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c
result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c
result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c
result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c
tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_cond,
tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_left,
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_right,
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3
tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_cond,
tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue,
tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse,
tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_left,
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_right,
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output,
 sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output,
 tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1525_c3_1635 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1529_c3_6da8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1535_c22_e01a_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1539_c22_b216_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1544_c3_f2c0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_2c93_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_94b6_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1531_l1523_l1528_DUPLICATE_106a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1531_l1537_l1541_DUPLICATE_4faf_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1552_l1519_DUPLICATE_2f80_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1544_c3_f2c0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1544_c3_f2c0;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1529_c3_6da8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1529_c3_6da8;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1525_c3_1635 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1525_c3_1635;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1541_c11_d466] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_left;
     BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output := BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1531_l1523_l1528_DUPLICATE_106a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1531_l1523_l1528_DUPLICATE_106a_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1539_c22_b216] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1539_c22_b216_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1537_c11_8e86] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_left;
     BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output := BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1534_c30_60ef] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_ins;
     sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_x;
     sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output := sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1531_l1537_l1541_DUPLICATE_4faf LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1531_l1537_l1541_DUPLICATE_4faf_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1528_c11_7086] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_left;
     BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output := BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1547_c11_8f7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1531_c11_f311] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_left;
     BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output := BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_2c93 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_2c93_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1523_c6_295a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1535_c22_e01a] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1535_c22_e01a_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_94b6 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_94b6_return_output := result.u16_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c6_295a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1528_c11_7086_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1531_c11_f311_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1537_c11_8e86_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_d466_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_8f7e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1535_c22_e01a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1539_c22_b216_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1531_l1523_l1528_DUPLICATE_106a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1531_l1523_l1528_DUPLICATE_106a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1531_l1523_l1528_DUPLICATE_106a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_94b6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_94b6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_94b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1547_l1541_l1537_l1531_l1528_DUPLICATE_1fe5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_2c93_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_2c93_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1523_l1537_l1528_DUPLICATE_2c93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1523_l1547_l1537_l1531_l1528_DUPLICATE_8cc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1531_l1537_l1541_DUPLICATE_4faf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1531_l1537_l1541_DUPLICATE_4faf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1531_l1537_l1541_DUPLICATE_4faf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1523_l1541_l1537_l1531_l1528_DUPLICATE_7d5d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1534_c30_60ef_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1523_c1_0ab8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1541_c7_94b3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1547_c7_cd18] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1541_c7_94b3] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_cond;
     tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output := tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1547_c7_cd18] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1541_c7_94b3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1523_c1_0ab8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_cd18_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;
     -- printf_uxn_opcodes_h_l1524_c3_43be[uxn_opcodes_h_l1524_c3_43be] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1524_c3_43be_uxn_opcodes_h_l1524_c3_43be_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u16_value_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1541_c7_94b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     t8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     t8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1541_c7_94b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_94b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- t8_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     t8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     t8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1537_c7_b42c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1537_c7_b42c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1531_c7_5c81] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1531_c7_5c81_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1528_c7_9392] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1528_c7_9392_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1523_c2_f166] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1552_l1519_DUPLICATE_2f80 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1552_l1519_DUPLICATE_2f80_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_284d(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c2_f166_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c2_f166_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1552_l1519_DUPLICATE_2f80_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1552_l1519_DUPLICATE_2f80_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
