-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity ldr_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_f74745d5;
architecture arch of ldr_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1622_c6_b60a]
signal BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1622_c2_6ca4]
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1635_c11_8bb0]
signal BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1635_c7_436c]
signal t8_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1635_c7_436c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1635_c7_436c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1635_c7_436c]
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1635_c7_436c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1635_c7_436c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1635_c7_436c]
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1635_c7_436c]
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1638_c11_6885]
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1638_c7_d468]
signal t8_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1638_c7_d468]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1638_c7_d468]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1638_c7_d468]
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1638_c7_d468]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1638_c7_d468]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1638_c7_d468]
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1638_c7_d468]
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1640_c30_e041]
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1641_c22_09c5]
signal BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1643_c11_849b]
signal BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1643_c7_10ca]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1643_c7_10ca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1643_c7_10ca]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1643_c7_10ca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1643_c7_10ca]
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1643_c7_10ca]
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1646_c11_422f]
signal BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1646_c7_ebd0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1646_c7_ebd0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1646_c7_ebd0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1646_c7_ebd0]
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1646_c7_ebd0]
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(7 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_left,
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_right,
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output);

-- t8_MUX_uxn_opcodes_h_l1622_c2_6ca4
t8_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4
tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond,
tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue,
tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse,
tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_left,
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_right,
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output);

-- t8_MUX_uxn_opcodes_h_l1635_c7_436c
t8_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
t8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
t8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1635_c7_436c
tmp8_MUX_uxn_opcodes_h_l1635_c7_436c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_cond,
tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_left,
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_right,
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output);

-- t8_MUX_uxn_opcodes_h_l1638_c7_d468
t8_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
t8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
t8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1638_c7_d468
tmp8_MUX_uxn_opcodes_h_l1638_c7_d468 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_cond,
tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue,
tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse,
tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1640_c30_e041
sp_relative_shift_uxn_opcodes_h_l1640_c30_e041 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_ins,
sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_x,
sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_y,
sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_left,
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_right,
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_left,
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_right,
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_cond,
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca
tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_cond,
tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue,
tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse,
tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_left,
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_right,
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0
tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond,
tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue,
tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse,
tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output,
 t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output,
 t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output,
 t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output,
 sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output,
 tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output,
 tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1627_c3_827f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1632_c3_5d2f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1636_c3_f2ab : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1641_c3_74d9 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1641_c27_e4a4_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1644_c3_6cc3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1649_c3_7745 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1622_l1635_l1638_DUPLICATE_2b30_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1643_l1635_DUPLICATE_f20e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1643_l1646_l1638_DUPLICATE_5047_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1654_l1618_DUPLICATE_3fb2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1636_c3_f2ab := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1636_c3_f2ab;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1627_c3_827f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1627_c3_827f;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1649_c3_7745 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1649_c3_7745;
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1632_c3_5d2f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1632_c3_5d2f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1644_c3_6cc3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1644_c3_6cc3;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse := tmp8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1622_l1635_l1638_DUPLICATE_2b30 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1622_l1635_l1638_DUPLICATE_2b30_return_output := result.u16_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1622_c6_b60a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1635_c11_8bb0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1643_l1635_DUPLICATE_f20e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1643_l1635_DUPLICATE_f20e_return_output := result.sp_relative_shift;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1641_c27_e4a4] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1641_c27_e4a4_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1643_c11_849b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1643_l1646_l1638_DUPLICATE_5047 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1643_l1646_l1638_DUPLICATE_5047_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1646_c11_422f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1640_c30_e041] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_ins;
     sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_x;
     sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output := sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1638_c11_6885] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_left;
     BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output := BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_b60a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_8bb0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_6885_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_849b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_422f_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1641_c27_e4a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1643_l1635_DUPLICATE_f20e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1643_l1635_DUPLICATE_f20e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1622_l1635_l1638_DUPLICATE_2b30_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1622_l1635_l1638_DUPLICATE_2b30_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1622_l1635_l1638_DUPLICATE_2b30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_0a4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1643_l1635_l1646_l1638_DUPLICATE_9c96_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1643_l1646_l1638_DUPLICATE_5047_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1643_l1646_l1638_DUPLICATE_5047_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1643_l1646_l1638_DUPLICATE_5047_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1622_l1646_l1643_l1638_l1635_DUPLICATE_77aa_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1622_c2_6ca4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_e041_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1643_c7_10ca] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1646_c7_ebd0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1646_c7_ebd0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     t8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     t8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1641_c22_09c5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1646_c7_ebd0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond;
     tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output := tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1646_c7_ebd0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1646_c7_ebd0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1641_c3_74d9 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_09c5_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_ebd0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1641_c3_74d9;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1643_c7_10ca] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1643_c7_10ca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1643_c7_10ca] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output := result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1643_c7_10ca] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_cond;
     tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output := tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1643_c7_10ca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- t8_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     t8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     t8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_10ca_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1638_c7_d468] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_cond;
     tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output := tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_d468_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1635_c7_436c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_436c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1622_c2_6ca4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1654_l1618_DUPLICATE_3fb2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1654_l1618_DUPLICATE_3fb2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_6ca4_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1654_l1618_DUPLICATE_3fb2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1654_l1618_DUPLICATE_3fb2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
