-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity nip_0CLK_6481cb28 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip_0CLK_6481cb28;
architecture arch of nip_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1870_c6_a832]
signal BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1870_c1_e4f9]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal t8_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1870_c2_89e1]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1871_c3_0129[uxn_opcodes_h_l1871_c3_0129]
signal printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1876_c11_6516]
signal BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1876_c7_0f1f]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1879_c11_9009]
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal t8_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1879_c7_0f72]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1883_c32_f26d]
signal BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1883_c32_de36]
signal BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1883_c32_dbb0]
signal MUX_uxn_opcodes_h_l1883_c32_dbb0_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1883_c32_dbb0_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1883_c32_dbb0_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1885_c11_2122]
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1885_c7_9a45]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1885_c7_9a45]
signal result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1885_c7_9a45]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1885_c7_9a45]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1885_c7_9a45]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1891_c11_02eb]
signal BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1891_c7_db3e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1891_c7_db3e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e56b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_stack_read := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832
BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_left,
BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_right,
BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output);

-- t8_MUX_uxn_opcodes_h_l1870_c2_89e1
t8_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1
result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1
result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1
result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1
result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1
result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

-- printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129
printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129 : entity work.printf_uxn_opcodes_h_l1871_c3_0129_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516
BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_left,
BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_right,
BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output);

-- t8_MUX_uxn_opcodes_h_l1876_c7_0f1f
t8_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f
result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_left,
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_right,
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output);

-- t8_MUX_uxn_opcodes_h_l1879_c7_0f72
t8_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72
result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72
result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d
BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_left,
BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_right,
BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36
BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_left,
BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_right,
BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output);

-- MUX_uxn_opcodes_h_l1883_c32_dbb0
MUX_uxn_opcodes_h_l1883_c32_dbb0 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1883_c32_dbb0_cond,
MUX_uxn_opcodes_h_l1883_c32_dbb0_iftrue,
MUX_uxn_opcodes_h_l1883_c32_dbb0_iffalse,
MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_left,
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_right,
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45
result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_cond,
result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb
BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_left,
BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_right,
BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e
result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e
result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output,
 t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output,
 t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output,
 t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output,
 MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1873_c3_fb8d : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1877_c3_3b37 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1888_c3_4dce : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1870_l1885_l1876_DUPLICATE_657b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1879_l1870_l1876_DUPLICATE_da3d_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1879_l1876_DUPLICATE_76ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1879_l1885_DUPLICATE_4d27_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1896_l1866_DUPLICATE_9e3b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_right := to_unsigned(128, 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1873_c3_fb8d := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1873_c3_fb8d;
     VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_iffalse := resize(to_signed(-1, 2), 8);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_right := to_unsigned(3, 2);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1877_c3_3b37 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1877_c3_3b37;
     VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1888_c3_4dce := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1888_c3_4dce;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1870_c6_a832] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_left;
     BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output := BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1870_l1885_l1876_DUPLICATE_657b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1870_l1885_l1876_DUPLICATE_657b_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1879_l1876_DUPLICATE_76ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1879_l1876_DUPLICATE_76ba_return_output := result.is_stack_read;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911_return_output := result.is_stack_write;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1879_l1870_l1876_DUPLICATE_da3d LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1879_l1870_l1876_DUPLICATE_da3d_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1891_c11_02eb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1879_l1885_DUPLICATE_4d27 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1879_l1885_DUPLICATE_4d27_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0_return_output := result.stack_value;

     -- BIN_OP_AND[uxn_opcodes_h_l1883_c32_f26d] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_left;
     BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output := BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1885_c11_2122] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_left;
     BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output := BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1876_c11_6516] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_left;
     BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output := BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1879_c11_9009] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_left;
     BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output := BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1883_c32_f26d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1870_c6_a832_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1876_c11_6516_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_9009_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_2122_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1891_c11_02eb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1879_l1870_l1876_DUPLICATE_da3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1879_l1870_l1876_DUPLICATE_da3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1879_l1870_l1876_DUPLICATE_da3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1879_l1885_l1876_l1891_DUPLICATE_3082_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1870_l1885_l1876_DUPLICATE_657b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1870_l1885_l1876_DUPLICATE_657b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1870_l1885_l1876_DUPLICATE_657b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1879_l1876_DUPLICATE_76ba_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1879_l1876_DUPLICATE_76ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1879_l1870_l1876_l1891_DUPLICATE_0911_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1879_l1885_DUPLICATE_4d27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1879_l1885_DUPLICATE_4d27_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1879_l1870_l1885_l1876_DUPLICATE_e7f0_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1885_c7_9a45] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1891_c7_db3e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1870_c1_e4f9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1891_c7_db3e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1885_c7_9a45] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output := result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;

     -- t8_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1883_c32_de36] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_left;
     BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output := BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1885_c7_9a45] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1883_c32_de36_return_output;
     VAR_printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1870_c1_e4f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1891_c7_db3e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1885_c7_9a45] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;

     -- MUX[uxn_opcodes_h_l1883_c32_dbb0] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1883_c32_dbb0_cond <= VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_cond;
     MUX_uxn_opcodes_h_l1883_c32_dbb0_iftrue <= VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_iftrue;
     MUX_uxn_opcodes_h_l1883_c32_dbb0_iffalse <= VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output := MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- printf_uxn_opcodes_h_l1871_c3_0129[uxn_opcodes_h_l1871_c3_0129] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1871_c3_0129_uxn_opcodes_h_l1871_c3_0129_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- t8_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1885_c7_9a45] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue := VAR_MUX_uxn_opcodes_h_l1883_c32_dbb0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_9a45_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     -- result_is_stack_read_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1879_c7_0f72] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;

     -- t8_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_0f72_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1876_c7_0f1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1876_c7_0f1f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1870_c2_89e1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1896_l1866_DUPLICATE_9e3b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1896_l1866_DUPLICATE_9e3b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e56b(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1870_c2_89e1_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1896_l1866_DUPLICATE_9e3b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1896_l1866_DUPLICATE_9e3b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
