-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_bce25fe8;
architecture arch of sta_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2299_c6_ebb3]
signal BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal t16_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal n8_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2299_c2_8a15]
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2312_c11_31aa]
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal t16_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal n8_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2312_c7_caa1]
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_8897]
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_3b1f]
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2317_c3_fcec]
signal CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2320_c11_77c6]
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal t16_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal n8_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2320_c7_be0c]
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2321_c3_8184]
signal BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_3dbf]
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2323_c7_e61a]
signal n8_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2323_c7_e61a]
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_e61a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_e61a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2323_c7_e61a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_e61a]
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2325_c30_8ff6]
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a906( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.u8_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_left,
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_right,
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output);

-- t16_MUX_uxn_opcodes_h_l2299_c2_8a15
t16_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- n8_MUX_uxn_opcodes_h_l2299_c2_8a15
n8_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond,
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_left,
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_right,
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output);

-- t16_MUX_uxn_opcodes_h_l2312_c7_caa1
t16_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- n8_MUX_uxn_opcodes_h_l2312_c7_caa1
n8_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_left,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_right,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output);

-- t16_MUX_uxn_opcodes_h_l2315_c7_3b1f
t16_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- n8_MUX_uxn_opcodes_h_l2315_c7_3b1f
n8_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec
CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_x,
CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_left,
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_right,
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output);

-- t16_MUX_uxn_opcodes_h_l2320_c7_be0c
t16_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- n8_MUX_uxn_opcodes_h_l2320_c7_be0c
n8_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184
BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_left,
BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_right,
BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_left,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_right,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output);

-- n8_MUX_uxn_opcodes_h_l2323_c7_e61a
n8_MUX_uxn_opcodes_h_l2323_c7_e61a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2323_c7_e61a_cond,
n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue,
n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse,
n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond,
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6
sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_ins,
sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_x,
sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_y,
sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output,
 t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output,
 t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output,
 t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output,
 CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output,
 t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output,
 n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output,
 sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_70dc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2304_c3_7505 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_eb1b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_3339 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2315_c7_3b1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2321_l2316_DUPLICATE_70cf_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l2332_l2294_DUPLICATE_b5dc_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_70dc := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_70dc;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_3339 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_3339;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_eb1b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_eb1b;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2304_c3_7505 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2304_c3_7505;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := t16;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_3dbf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output := result.u8_value;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output := result.is_stack_write;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2321_l2316_DUPLICATE_70cf LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2321_l2316_DUPLICATE_70cf_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2312_c11_31aa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2320_c11_77c6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2325_c30_8ff6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_ins;
     sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_x;
     sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output := sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output := result.u16_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2315_c7_3b1f_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2299_c6_ebb3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_8897] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_left;
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output := BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_ebb3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_31aa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_8897_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_77c6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_3dbf_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2321_l2316_DUPLICATE_70cf_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2321_l2316_DUPLICATE_70cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_ded4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_8005_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_13dd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2320_l2312_l2323_l2315_DUPLICATE_d3bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2312_l2299_l2323_l2320_l2315_DUPLICATE_6873_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2299_c2_8a15_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_8ff6_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2321_c3_8184] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_left;
     BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output := BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_e61a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_e61a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_e61a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- n8_MUX[uxn_opcodes_h_l2323_c7_e61a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2323_c7_e61a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_cond;
     n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue;
     n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output := n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2317_c3_fcec] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output := CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2323_c7_e61a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2323_c7_e61a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output := result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_8184_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_fcec_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_e61a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- t16_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2320_c7_be0c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2320_c7_be0c_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- t16_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c7_3b1f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2315_c7_3b1f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- n8_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- t16_MUX[uxn_opcodes_h_l2312_c7_caa1] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2312_c7_caa1_cond <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_cond;
     t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iftrue;
     t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output := t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2312_c7_caa1_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- t16_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- n8_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2299_c2_8a15] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output := result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l2332_l2294_DUPLICATE_b5dc LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l2332_l2294_DUPLICATE_b5dc_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a906(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_8a15_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l2332_l2294_DUPLICATE_b5dc_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l2332_l2294_DUPLICATE_b5dc_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
