-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2236_c6_47e2]
signal BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2236_c2_3b3a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2249_c11_d754]
signal BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2249_c7_1002]
signal t8_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2249_c7_1002]
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2249_c7_1002]
signal n8_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2249_c7_1002]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2249_c7_1002]
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2249_c7_1002]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2249_c7_1002]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2249_c7_1002]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2252_c11_519b]
signal BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2252_c7_c4d0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2254_c30_b55e]
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2256_c11_3b20]
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2256_c7_e329]
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2256_c7_e329]
signal n8_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2256_c7_e329]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2256_c7_e329]
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2256_c7_e329]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2256_c7_e329]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2256_c7_e329]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2259_c18_1656]
signal BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2259_c11_41ca]
signal BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2259_c34_c6ed]
signal CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2259_c11_9b26]
signal BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_left,
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_right,
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output);

-- t8_MUX_uxn_opcodes_h_l2236_c2_3b3a
t8_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a
tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- n8_MUX_uxn_opcodes_h_l2236_c2_3b3a
n8_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_left,
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_right,
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output);

-- t8_MUX_uxn_opcodes_h_l2249_c7_1002
t8_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
t8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
t8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2249_c7_1002
tmp8_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- n8_MUX_uxn_opcodes_h_l2249_c7_1002
n8_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
n8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
n8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_left,
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_right,
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output);

-- t8_MUX_uxn_opcodes_h_l2252_c7_c4d0
t8_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0
tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- n8_MUX_uxn_opcodes_h_l2252_c7_c4d0
n8_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e
sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_ins,
sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_x,
sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_y,
sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_left,
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_right,
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2256_c7_e329
tmp8_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- n8_MUX_uxn_opcodes_h_l2256_c7_e329
n8_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
n8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
n8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656
BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_left,
BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_right,
BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca
BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_left,
BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_right,
BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed
CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_x,
CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26
BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26 : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_left,
BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_right,
BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output,
 t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output,
 t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output,
 t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output,
 sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output,
 tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output,
 CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2241_c3_6b7f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2246_c3_cc19 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2250_c3_b556 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2258_c3_f381 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_cbc3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_e3f1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_c2dc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_2335_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2256_l2252_DUPLICATE_f8d0_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2266_l2232_DUPLICATE_6db0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_cbc3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_cbc3;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2258_c3_f381 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2258_c3_f381;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2241_c3_6b7f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2241_c3_6b7f;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2250_c3_b556 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2250_c3_b556;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_right := to_unsigned(15, 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2246_c3_cc19 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2246_c3_cc19;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := tmp8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_c2dc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_c2dc_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output := result.is_stack_index_flipped;

     -- CONST_SR_4[uxn_opcodes_h_l2259_c34_c6ed] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output := CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_e3f1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_e3f1_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2249_c11_d754] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_left;
     BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output := BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2252_c11_519b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2254_c30_b55e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_ins;
     sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_x;
     sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output := sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2236_c6_47e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2256_l2252_DUPLICATE_f8d0 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2256_l2252_DUPLICATE_f8d0_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_2335 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_2335_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2256_c11_3b20] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_left;
     BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output := BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2259_c18_1656] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_left;
     BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output := BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_1656_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_47e2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_d754_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_519b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_3b20_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_c2dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_c2dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_e3f1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_e3f1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_e3f1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_2335_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_2335_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2256_l2249_l2252_DUPLICATE_2335_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2256_l2252_DUPLICATE_f8d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2256_l2252_DUPLICATE_f8d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2236_l2256_l2249_l2252_DUPLICATE_3b2c_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_right := VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_c6ed_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_b55e_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2259_c11_41ca] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_left;
     BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output := BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- n8_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     n8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     n8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- t8_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_41ca_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     t8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     t8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- n8_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2259_c11_9b26] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_left;
     BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output := BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_9b26_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     -- t8_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2256_c7_e329] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output := result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;

     -- n8_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     n8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     n8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e329_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2252_c7_c4d0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c4d0_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2249_c7_1002] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output := result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1002_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2236_c2_3b3a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_cond;
     tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output := tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2266_l2232_DUPLICATE_6db0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2266_l2232_DUPLICATE_6db0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_3b3a_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2266_l2232_DUPLICATE_6db0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2266_l2232_DUPLICATE_6db0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
