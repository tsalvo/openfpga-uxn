-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_16;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint8_t_array_16_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iftrue : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iffalse : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iftrue : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iffalse : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iftrue : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iffalse : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iftrue : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iffalse : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iftrue : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iffalse : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iftrue : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iffalse : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iftrue : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iffalse : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iftrue : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iffalse : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_f08f( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_array_16_t is
 
  variable base : uint8_t_array_16_t; 
  variable return_output : uint8_t_array_16_t;
begin
      base.data(0) := ref_toks_0;
      base.data(3) := ref_toks_1;
      base.data(9) := ref_toks_2;
      base.data(6) := ref_toks_3;
      base.data(12) := ref_toks_4;
      base.data(15) := ref_toks_5;
      base.data(4) := ref_toks_6;
      base.data(1) := ref_toks_7;
      base.data(7) := ref_toks_8;
      base.data(10) := ref_toks_9;
      base.data(13) := ref_toks_10;
      base.data(2) := ref_toks_11;
      base.data(5) := ref_toks_12;
      base.data(8) := ref_toks_13;
      base.data(14) := ref_toks_14;
      base.data(11) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_16;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint8_t_array_16_t;
 variable VAR_base : uint8_t_16;
 variable VAR_rv : uint8_t_array_16_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_0ad2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_2593_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_28ba_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c15_7642_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_f414_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_ce0d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_b6ca_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_99b4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_30dc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_eee9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4f39_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_ed12_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8b65_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_aad4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_e1b2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_e8e1_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_f08f_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0059_return_output : uint8_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_right := to_unsigned(14, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_12_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_f414] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_f414_return_output := VAR_ref_toks_0(12);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_2593] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_2593_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_16_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_ed12] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_ed12_return_output := VAR_ref_toks_0(2);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_99b4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_99b4_return_output := VAR_ref_toks_0(1);

     -- CONST_REF_RD_uint8_t_uint8_t_16_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8b65] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8b65_return_output := VAR_ref_toks_0(5);

     -- CONST_REF_RD_uint8_t_uint8_t_16_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c15_7642] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c15_7642_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_16_13_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4f39] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4f39_return_output := VAR_ref_toks_0(13);

     -- CONST_REF_RD_uint8_t_uint8_t_16_14_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_e1b2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_e1b2_return_output := VAR_ref_toks_0(14);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_30dc] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_30dc_return_output := VAR_ref_toks_0(7);

     -- CONST_REF_RD_uint8_t_uint8_t_16_8_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_aad4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_aad4_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_16_15_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_ce0d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_ce0d_return_output := VAR_ref_toks_0(15);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_0ad2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_0ad2_return_output := VAR_ref_toks_0(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_10_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_eee9] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_eee9_return_output := VAR_ref_toks_0(10);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_9_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_28ba] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_28ba_return_output := VAR_ref_toks_0(9);

     -- CONST_REF_RD_uint8_t_uint8_t_16_11_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_e8e1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_e8e1_return_output := VAR_ref_toks_0(11);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_b6ca] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_b6ca_return_output := VAR_ref_toks_0(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output;

     -- Submodule level 1
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_5161_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_e074_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_d5e5_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3f89_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d330_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_df41_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ef66_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_be84_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_52b4_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_06f2_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_bc39_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_bfa5_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_3d20_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_68dd_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_2420_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_7f0a_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_0ad2_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_eee9_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_e8e1_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_f414_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4f39_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_e1b2_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_ce0d_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_99b4_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_ed12_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_2593_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_b6ca_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8b65_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c15_7642_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_30dc_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_aad4_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_28ba_return_output;
     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322] LATENCY=0
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_iffalse;
     -- Outputs
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c] LATENCY=0
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_iffalse;
     -- Outputs
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679] LATENCY=0
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_iffalse;
     -- Outputs
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5] LATENCY=0
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_iffalse;
     -- Outputs
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906] LATENCY=0
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_iffalse;
     -- Outputs
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11] LATENCY=0
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_iffalse;
     -- Outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b] LATENCY=0
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_iffalse;
     -- Outputs
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08] LATENCY=0
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_iffalse;
     -- Outputs
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_f08f[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0059] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_f08f_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0059_return_output := CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_f08f(
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_09e1_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_e8b3_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_c679_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_245f_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_f906_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b43c_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_ae38_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_4c3c_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7c34_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_7c11_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_2322_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_5051_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_080d_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_ba08_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_e4b5_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_9a3b_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_f08f_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0059_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
