-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity sft2_0CLK_91f0cf2d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end sft2_0CLK_91f0cf2d;
architecture arch of sft2_0CLK_91f0cf2d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2032_c6_08d1]
signal BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(7 downto 0);

-- n16_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2032_c2_0eb5]
signal tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2039_c11_3910]
signal BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal t8_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(7 downto 0);

-- n16_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal n16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2039_c7_ae82]
signal tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2043_c11_a2b2]
signal BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2043_c7_8486]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2043_c7_8486]
signal t8_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(7 downto 0);

-- n16_MUX[uxn_opcodes_h_l2043_c7_8486]
signal n16_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2043_c7_8486]
signal tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2046_c30_7ff6]
signal sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2048_c11_7dfe]
signal BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2048_c7_e630]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2048_c7_e630]
signal result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2048_c7_e630]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2048_c7_e630]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2048_c7_e630]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2048_c7_e630]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l2048_c7_e630]
signal n16_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2048_c7_e630]
signal tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(15 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2050_c20_6882]
signal BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2050_c12_9ed1]
signal BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_left : unsigned(15 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output : unsigned(15 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2050_c36_ca3e]
signal CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2050_c12_0f1c]
signal BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_left : unsigned(15 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2056_c11_9965]
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2056_c7_ebd4]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c7_ebd4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c7_ebd4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1
BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_left,
BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_right,
BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- t8_MUX_uxn_opcodes_h_l2032_c2_0eb5
t8_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- n16_MUX_uxn_opcodes_h_l2032_c2_0eb5
n16_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5
tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond,
tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue,
tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse,
tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910
BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_left,
BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_right,
BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82
result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82
result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82
result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82
result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82
result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- t8_MUX_uxn_opcodes_h_l2039_c7_ae82
t8_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- n16_MUX_uxn_opcodes_h_l2039_c7_ae82
n16_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82
tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond,
tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue,
tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse,
tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2
BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_left,
BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_right,
BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486
result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486
result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486
result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486
result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486
result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- t8_MUX_uxn_opcodes_h_l2043_c7_8486
t8_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
t8_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
t8_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- n16_MUX_uxn_opcodes_h_l2043_c7_8486
n16_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
n16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
n16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2043_c7_8486
tmp16_MUX_uxn_opcodes_h_l2043_c7_8486 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_cond,
tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue,
tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse,
tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6
sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_ins,
sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_x,
sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_y,
sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe
BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_left,
BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_right,
BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630
result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630
result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630
result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630
result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- n16_MUX_uxn_opcodes_h_l2048_c7_e630
n16_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
n16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
n16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2048_c7_e630
tmp16_MUX_uxn_opcodes_h_l2048_c7_e630 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_cond,
tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue,
tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse,
tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882
BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_left,
BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_right,
BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1
BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1 : entity work.BIN_OP_SR_uint16_t_uint8_t_0CLK_295015b8 port map (
BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_left,
BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_right,
BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e
CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_x,
CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c
BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c : entity work.BIN_OP_SL_uint16_t_uint8_t_0CLK_b6546dec port map (
BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_left,
BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_right,
BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965
BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_left,
BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_right,
BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output,
 sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output,
 CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2036_c3_5e6f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2041_c3_be33 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2044_c8_5730_return_output : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2053_c3_80f9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2032_l2048_l2039_DUPLICATE_4432_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2043_l2032_l2039_DUPLICATE_df61_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2043_l2048_DUPLICATE_c910_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2062_l2027_DUPLICATE_67cc_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_right := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_right := to_unsigned(15, 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2053_c3_80f9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2053_c3_80f9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_right := to_unsigned(3, 2);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2041_c3_be33 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2041_c3_be33;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2036_c3_5e6f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2036_c3_5e6f;
     VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := t8;
     VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2056_c11_9965] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_left;
     BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output := BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2046_c30_7ff6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_ins;
     sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_x;
     sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output := sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2043_l2032_l2039_DUPLICATE_df61 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2043_l2032_l2039_DUPLICATE_df61_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2048_c11_7dfe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_left;
     BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output := BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2032_c6_08d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2050_c20_6882] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_left;
     BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output := BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2032_l2048_l2039_DUPLICATE_4432 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2032_l2048_l2039_DUPLICATE_4432_return_output := result.is_sp_shift;

     -- CONST_SR_4[uxn_opcodes_h_l2050_c36_ca3e] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output := CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2044_c8_5730] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2044_c8_5730_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2039_c11_3910] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_left;
     BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output := BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62_return_output := result.u16_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2043_l2048_DUPLICATE_c910 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2043_l2048_DUPLICATE_c910_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2043_c11_a2b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7_return_output := result.is_stack_operation_16bit;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2050_c20_6882_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c6_08d1_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2039_c11_3910_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2043_c11_a2b2_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2048_c11_7dfe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c11_9965_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2044_c8_5730_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2043_l2032_l2039_DUPLICATE_df61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2043_l2032_l2039_DUPLICATE_df61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2043_l2032_l2039_DUPLICATE_df61_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2039_DUPLICATE_4d62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2043_l2048_l2039_l2056_DUPLICATE_a9f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2032_l2048_l2039_DUPLICATE_4432_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2032_l2048_l2039_DUPLICATE_4432_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2032_l2048_l2039_DUPLICATE_4432_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2043_l2032_l2048_l2056_DUPLICATE_34e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2043_l2032_l2039_l2056_DUPLICATE_82eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2043_l2048_DUPLICATE_c910_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2043_l2048_DUPLICATE_c910_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_right := VAR_CONST_SR_4_uxn_opcodes_h_l2050_c36_ca3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2046_c30_7ff6_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2056_c7_ebd4] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c7_ebd4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c7_ebd4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- t8_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     t8_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     t8_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2050_c12_9ed1] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_left;
     BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output := BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output;

     -- n16_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     n16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     n16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2050_c12_9ed1_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c7_ebd4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- t8_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- n16_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     n16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     n16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2050_c12_0f1c] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_left;
     BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output := BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- Submodule level 3
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2050_c12_0f1c_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     -- n16_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- t8_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2048_c7_e630] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_cond;
     tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output := tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2048_c7_e630_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2043_c7_8486] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_cond;
     tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output := tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;

     -- n16_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2043_c7_8486_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2039_c7_ae82] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output := result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;

     -- Submodule level 6
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2039_c7_ae82_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2032_c2_0eb5] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_cond;
     tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output := tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;

     -- Submodule level 7
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2062_l2027_DUPLICATE_67cc LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2062_l2027_DUPLICATE_67cc_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c2_0eb5_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2062_l2027_DUPLICATE_67cc_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2062_l2027_DUPLICATE_67cc_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
