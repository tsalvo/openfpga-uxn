-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_8167]
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2419_c2_2be3]
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_7949]
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2432_c7_6298]
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_6298]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_6298]
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_6298]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_6298]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_6298]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_6298]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2432_c7_6298]
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_ed22]
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2435_c7_a793]
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_a793]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_a793]
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_a793]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_a793]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_a793]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_a793]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2435_c7_a793]
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2437_c30_e8d1]
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_1333]
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_2eee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_9e05]
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_2c8a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_2c8a]
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_2c8a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_2c8a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_left,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_right,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3
t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3
t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_cond,
t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue,
t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse,
t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_left,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_right,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2432_c7_6298
t16_low_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2432_c7_6298
t16_high_MUX_uxn_opcodes_h_l2432_c7_6298 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_cond,
t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue,
t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse,
t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_left,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_right,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2435_c7_a793
t16_low_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2435_c7_a793
t16_high_MUX_uxn_opcodes_h_l2435_c7_a793 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_cond,
t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue,
t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse,
t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1
sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_ins,
sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_x,
sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_y,
sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_left,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_right,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee
t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_left,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_right,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output,
 t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output,
 t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output,
 t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output,
 sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output,
 t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_32b5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_1a55 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_b861 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_594a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_4fe2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_f7d6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_1cd7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_a14c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_dbda_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_ae89_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2435_l2447_DUPLICATE_6195_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2415_l2454_DUPLICATE_8c1e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_b861 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_b861;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_f7d6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_f7d6;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_4fe2 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_4fe2;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_32b5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_32b5;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_1a55 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_1a55;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_1cd7 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_1cd7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_594a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_594a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_right := to_unsigned(4, 3);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_y := resize(to_signed(-2, 3), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_9e05] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_left;
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output := BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_ed22] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_left;
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output := BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_1333] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_left;
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output := BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_a14c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_a14c_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_8167] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_left;
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output := BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_dbda LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_dbda_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2437_c30_e8d1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_ins;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_x;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output := sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_7949] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_left;
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output := BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2435_l2447_DUPLICATE_6195 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2435_l2447_DUPLICATE_6195_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_ae89 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_ae89_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_8167_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7949_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_ed22_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_1333_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_9e05_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_ae89_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_ae89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2435_l2439_l2432_l2447_DUPLICATE_7e6f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_a14c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_a14c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_a14c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_dbda_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_dbda_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2435_l2439_l2432_DUPLICATE_dbda_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2435_l2447_DUPLICATE_6195_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2435_l2447_DUPLICATE_6195_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2435_l2419_l2432_l2447_DUPLICATE_4219_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_2be3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_e8d1_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_2c8a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_2c8a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_2c8a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_2c8a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_2c8a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_2eee] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output := result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2eee_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_a793] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output := result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_a793_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_6298] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_6298_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_2be3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2415_l2454_DUPLICATE_8c1e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2415_l2454_DUPLICATE_8c1e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_2be3_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2415_l2454_DUPLICATE_8c1e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2415_l2454_DUPLICATE_8c1e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
