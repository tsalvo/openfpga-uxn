-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity nip_0CLK_4351dde2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip_0CLK_4351dde2;
architecture arch of nip_0CLK_4351dde2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1340_c6_e093]
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1340_c1_9914]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : signed(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1340_c2_bbc8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1341_c3_ce32[uxn_opcodes_h_l1341_c3_ce32]
signal printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1348_c11_26c6]
signal BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal t8_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : signed(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1348_c7_08d5]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1352_c11_7021]
signal BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1352_c7_5118]
signal t8_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : signed(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1352_c7_5118]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1356_c32_e22e]
signal BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1356_c32_b0ce]
signal BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1356_c32_0441]
signal MUX_uxn_opcodes_h_l1356_c32_0441_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1356_c32_0441_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1356_c32_0441_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1356_c32_0441_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1358_c11_db1b]
signal BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1358_c7_ab2e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1358_c7_ab2e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1358_c7_ab2e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1358_c7_ab2e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1358_c7_ab2e]
signal result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1364_c11_590a]
signal BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1364_c7_4f99]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1364_c7_4f99]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_49dd( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.stack_value := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_read := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_sp_shift := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093
BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_left,
BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_right,
BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output);

-- t8_MUX_uxn_opcodes_h_l1340_c2_bbc8
t8_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

-- printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32
printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32 : entity work.printf_uxn_opcodes_h_l1341_c3_ce32_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6
BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_left,
BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_right,
BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output);

-- t8_MUX_uxn_opcodes_h_l1348_c7_08d5
t8_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5
result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5
result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5
result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5
result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5
result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021
BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_left,
BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_right,
BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output);

-- t8_MUX_uxn_opcodes_h_l1352_c7_5118
t8_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
t8_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
t8_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118
result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118
result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118
result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118
result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118
result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118
result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e
BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_left,
BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_right,
BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce
BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_left,
BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_right,
BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output);

-- MUX_uxn_opcodes_h_l1356_c32_0441
MUX_uxn_opcodes_h_l1356_c32_0441 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1356_c32_0441_cond,
MUX_uxn_opcodes_h_l1356_c32_0441_iftrue,
MUX_uxn_opcodes_h_l1356_c32_0441_iffalse,
MUX_uxn_opcodes_h_l1356_c32_0441_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b
BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_left,
BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_right,
BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e
result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e
result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e
result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e
result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond,
result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a
BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_left,
BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_right,
BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99
result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99
result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output,
 t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output,
 t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output,
 t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output,
 MUX_uxn_opcodes_h_l1356_c32_0441_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1344_c3_080c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1350_c3_3c68 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1352_c7_5118_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1356_c32_0441_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1356_c32_0441_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1356_c32_0441_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1356_c32_0441_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1361_c3_e17c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1348_l1352_l1340_DUPLICATE_b5c2_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1348_l1358_l1340_DUPLICATE_7034_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1364_l1348_l1352_DUPLICATE_a5ad_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1358_l1352_DUPLICATE_357e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_49dd_uxn_opcodes_h_l1369_l1336_DUPLICATE_35ea_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_right := to_unsigned(128, 8);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1361_c3_e17c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1361_c3_e17c;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1356_c32_0441_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1344_c3_080c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1344_c3_080c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1350_c3_3c68 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1350_c3_3c68;
     VAR_MUX_uxn_opcodes_h_l1356_c32_0441_iffalse := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_right := to_unsigned(2, 2);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := t8;
     -- BIN_OP_AND[uxn_opcodes_h_l1356_c32_e22e] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_left;
     BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output := BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1340_c2_bbc8_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1364_l1348_l1352_DUPLICATE_a5ad LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1364_l1348_l1352_DUPLICATE_a5ad_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1348_c11_26c6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1352_c11_7021] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_left;
     BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output := BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1358_c11_db1b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1340_c6_e093] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_left;
     BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output := BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1348_l1358_l1340_DUPLICATE_7034 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1348_l1358_l1340_DUPLICATE_7034_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1358_l1352_DUPLICATE_357e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1358_l1352_DUPLICATE_357e_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1348_l1352_l1340_DUPLICATE_b5c2 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1348_l1352_l1340_DUPLICATE_b5c2_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1364_c11_590a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output;

     -- result_is_stack_read_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     VAR_result_is_stack_read_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1352_c7_5118_return_output := result.is_stack_read;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1356_c32_e22e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c6_e093_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1348_c11_26c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1352_c11_7021_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1358_c11_db1b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1364_c11_590a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1348_l1352_l1340_DUPLICATE_b5c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1348_l1352_l1340_DUPLICATE_b5c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1348_l1352_l1340_DUPLICATE_b5c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1364_DUPLICATE_6da5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1348_l1358_l1340_DUPLICATE_7034_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1348_l1358_l1340_DUPLICATE_7034_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1348_l1358_l1340_DUPLICATE_7034_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1364_l1348_l1352_DUPLICATE_a5ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1364_l1348_l1352_DUPLICATE_a5ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1364_l1348_l1352_DUPLICATE_a5ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1358_l1352_DUPLICATE_357e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1358_l1352_DUPLICATE_357e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1358_l1348_l1352_l1340_DUPLICATE_076e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1340_c2_bbc8_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_result_is_stack_read_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1352_c7_5118_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1364_c7_4f99] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1364_c7_4f99] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1356_c32_b0ce] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_left;
     BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output := BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1358_c7_ab2e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1358_c7_ab2e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1358_c7_ab2e] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output := result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1340_c1_9914] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     t8_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     t8_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1356_c32_0441_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1356_c32_b0ce_return_output;
     VAR_printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1340_c1_9914_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1364_c7_4f99_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     -- result_is_stack_read_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- t8_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1358_c7_ab2e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;

     -- MUX[uxn_opcodes_h_l1356_c32_0441] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1356_c32_0441_cond <= VAR_MUX_uxn_opcodes_h_l1356_c32_0441_cond;
     MUX_uxn_opcodes_h_l1356_c32_0441_iftrue <= VAR_MUX_uxn_opcodes_h_l1356_c32_0441_iftrue;
     MUX_uxn_opcodes_h_l1356_c32_0441_iffalse <= VAR_MUX_uxn_opcodes_h_l1356_c32_0441_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1356_c32_0441_return_output := MUX_uxn_opcodes_h_l1356_c32_0441_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1358_c7_ab2e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;

     -- printf_uxn_opcodes_h_l1341_c3_ce32[uxn_opcodes_h_l1341_c3_ce32] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1341_c3_ce32_uxn_opcodes_h_l1341_c3_ce32_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue := VAR_MUX_uxn_opcodes_h_l1356_c32_0441_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1358_c7_ab2e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- t8_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1352_c7_5118] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1352_c7_5118_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1348_c7_08d5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1348_c7_08d5_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1340_c2_bbc8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_49dd_uxn_opcodes_h_l1369_l1336_DUPLICATE_35ea LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_49dd_uxn_opcodes_h_l1369_l1336_DUPLICATE_35ea_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_49dd(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c2_bbc8_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_49dd_uxn_opcodes_h_l1369_l1336_DUPLICATE_35ea_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_49dd_uxn_opcodes_h_l1369_l1336_DUPLICATE_35ea_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
