-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity opc_neq_phased_0CLK_2ca51e56 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_neq_phased_0CLK_2ca51e56;
architecture arch of opc_neq_phased_0CLK_2ca51e56 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l448_c6_6dc8]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l448_c1_dffb]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l451_c7_39ed]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l448_c2_c7e2]
signal t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l448_c2_c7e2]
signal n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l448_c2_c7e2]
signal result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l449_c12_988e]
signal set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l451_c11_01dc]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l451_c1_9fc4]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l454_c7_3583]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l451_c7_39ed]
signal t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l451_c7_39ed]
signal n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l451_c7_39ed]
signal result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l452_c8_b4db]
signal t_register_uxn_opcodes_phased_h_l452_c8_b4db_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l454_c11_dfdd]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l454_c1_126b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l457_c7_324b]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l454_c7_3583]
signal t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l454_c7_3583]
signal n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l454_c7_3583]
signal result_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l455_c8_4786]
signal n_register_uxn_opcodes_phased_h_l455_c8_4786_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l457_c11_d9c2]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l457_c1_7500]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l460_c7_aab5]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l457_c7_324b]
signal n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l457_c7_324b]
signal result_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l458_c8_64e5]
signal n_register_uxn_opcodes_phased_h_l458_c8_64e5_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l460_c11_e8a3]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l460_c1_87fe]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l463_c7_2a27]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l460_c7_aab5]
signal result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l461_c3_f77d]
signal set_uxn_opcodes_phased_h_l461_c3_f77d_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l461_c3_f77d_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l461_c3_f77d_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l461_c3_f77d_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l461_c3_f77d_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l461_c3_f77d_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l461_c3_f77d_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l463_c11_2efa]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l463_c1_5b59]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l463_c7_2a27]
signal result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l464_c33_d30e]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_phased_h_l464_c33_b073]
signal MUX_uxn_opcodes_phased_h_l464_c33_b073_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_phased_h_l464_c33_b073_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_phased_h_l464_c33_b073_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_phased_h_l464_c3_4b11]
signal put_stack_uxn_opcodes_phased_h_l464_c3_4b11_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l464_c3_4b11_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l464_c3_4b11_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l464_c3_4b11_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l464_c3_4b11_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l466_c11_d282]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l466_c7_ae82]
signal result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8
BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2
t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond,
t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue,
t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse,
t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2
n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond,
n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue,
n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse,
n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output);

-- result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2
result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond,
result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue,
result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse,
result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l449_c12_988e
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_sp,
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_k,
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_mul,
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_add,
set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc
BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed
t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond,
t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue,
t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse,
t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed
n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond,
n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue,
n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse,
n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output);

-- result_MUX_uxn_opcodes_phased_h_l451_c7_39ed
result_MUX_uxn_opcodes_phased_h_l451_c7_39ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond,
result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue,
result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse,
result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output);

-- t_register_uxn_opcodes_phased_h_l452_c8_b4db
t_register_uxn_opcodes_phased_h_l452_c8_b4db : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l452_c8_b4db_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_index,
t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_ptr,
t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd
BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l454_c7_3583
t8_MUX_uxn_opcodes_phased_h_l454_c7_3583 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond,
t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue,
t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse,
t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l454_c7_3583
n8_MUX_uxn_opcodes_phased_h_l454_c7_3583 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond,
n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue,
n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse,
n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output);

-- result_MUX_uxn_opcodes_phased_h_l454_c7_3583
result_MUX_uxn_opcodes_phased_h_l454_c7_3583 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond,
result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue,
result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse,
result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output);

-- n_register_uxn_opcodes_phased_h_l455_c8_4786
n_register_uxn_opcodes_phased_h_l455_c8_4786 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l455_c8_4786_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_index,
n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_ptr,
n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2
BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l457_c7_324b
n8_MUX_uxn_opcodes_phased_h_l457_c7_324b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond,
n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue,
n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse,
n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output);

-- result_MUX_uxn_opcodes_phased_h_l457_c7_324b
result_MUX_uxn_opcodes_phased_h_l457_c7_324b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond,
result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue,
result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse,
result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output);

-- n_register_uxn_opcodes_phased_h_l458_c8_64e5
n_register_uxn_opcodes_phased_h_l458_c8_64e5 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l458_c8_64e5_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_index,
n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_ptr,
n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3
BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output);

-- result_MUX_uxn_opcodes_phased_h_l460_c7_aab5
result_MUX_uxn_opcodes_phased_h_l460_c7_aab5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond,
result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue,
result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse,
result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output);

-- set_uxn_opcodes_phased_h_l461_c3_f77d
set_uxn_opcodes_phased_h_l461_c3_f77d : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l461_c3_f77d_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l461_c3_f77d_sp,
set_uxn_opcodes_phased_h_l461_c3_f77d_stack_index,
set_uxn_opcodes_phased_h_l461_c3_f77d_ins,
set_uxn_opcodes_phased_h_l461_c3_f77d_k,
set_uxn_opcodes_phased_h_l461_c3_f77d_mul,
set_uxn_opcodes_phased_h_l461_c3_f77d_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa
BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output);

-- result_MUX_uxn_opcodes_phased_h_l463_c7_2a27
result_MUX_uxn_opcodes_phased_h_l463_c7_2a27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond,
result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue,
result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse,
result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e
BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output);

-- MUX_uxn_opcodes_phased_h_l464_c33_b073
MUX_uxn_opcodes_phased_h_l464_c33_b073 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_phased_h_l464_c33_b073_cond,
MUX_uxn_opcodes_phased_h_l464_c33_b073_iftrue,
MUX_uxn_opcodes_phased_h_l464_c33_b073_iffalse,
MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output);

-- put_stack_uxn_opcodes_phased_h_l464_c3_4b11
put_stack_uxn_opcodes_phased_h_l464_c3_4b11 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l464_c3_4b11_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l464_c3_4b11_sp,
put_stack_uxn_opcodes_phased_h_l464_c3_4b11_stack_index,
put_stack_uxn_opcodes_phased_h_l464_c3_4b11_offset,
put_stack_uxn_opcodes_phased_h_l464_c3_4b11_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282
BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output);

-- result_MUX_uxn_opcodes_phased_h_l466_c7_ae82
result_MUX_uxn_opcodes_phased_h_l466_c7_ae82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_cond,
result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iftrue,
result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iffalse,
result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output,
 t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output,
 n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output,
 result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output,
 set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output,
 t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output,
 n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output,
 result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output,
 t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output,
 t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output,
 n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output,
 result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output,
 n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output,
 n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output,
 result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output,
 n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output,
 result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output,
 result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output,
 MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output,
 result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_value : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_right := to_unsigned(5, 3);
     VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_add := resize(to_signed(-1, 2), 8);
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iffalse := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_offset := resize(to_unsigned(0, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_add := resize(to_signed(-1, 2), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_k := VAR_k;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_index := VAR_stack_index;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_right := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l464_c33_d30e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l448_c6_6dc8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l457_c11_d9c2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l466_c11_d282] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l454_c11_dfdd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l460_c11_e8a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l451_c11_01dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l463_c11_2efa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l448_c6_6dc8_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l451_c11_01dc_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l454_c11_dfdd_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l457_c11_d9c2_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l460_c11_e8a3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l463_c11_2efa_return_output;
     VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l464_c33_d30e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l466_c11_d282_return_output;
     -- MUX[uxn_opcodes_phased_h_l464_c33_b073] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_phased_h_l464_c33_b073_cond <= VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_cond;
     MUX_uxn_opcodes_phased_h_l464_c33_b073_iftrue <= VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_iftrue;
     MUX_uxn_opcodes_phased_h_l464_c33_b073_iffalse <= VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output := MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l466_c7_ae82] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_cond;
     result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iftrue;
     result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output := result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l451_c7_39ed] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l448_c1_dffb] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_value := VAR_MUX_uxn_opcodes_phased_h_l464_c33_b073_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l448_c1_dffb_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l466_c7_ae82_return_output;
     -- set_will_fail[uxn_opcodes_phased_h_l449_c12_988e] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_sp;
     set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_k;
     set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_mul;
     set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output := set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l451_c1_9fc4] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l463_c7_2a27] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond;
     result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue;
     result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output := result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l454_c7_3583] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l451_c1_9fc4_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l449_c12_988e_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l454_c1_126b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output;

     -- t_register[uxn_opcodes_phased_h_l452_c8_b4db] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l452_c8_b4db_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_index;
     t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output := t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l460_c7_aab5] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond;
     result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue;
     result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output := result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l457_c7_324b] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l454_c1_126b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue := VAR_t_register_uxn_opcodes_phased_h_l452_c8_b4db_return_output;
     -- n_register[uxn_opcodes_phased_h_l455_c8_4786] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l455_c8_4786_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_index;
     n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output := n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l457_c1_7500] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l457_c7_324b] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond;
     result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue;
     result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output := result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l460_c7_aab5] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c7_aab5_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l457_c1_7500_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue := VAR_n_register_uxn_opcodes_phased_h_l455_c8_4786_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l460_c1_87fe] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output;

     -- n_register[uxn_opcodes_phased_h_l458_c8_64e5] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l458_c8_64e5_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_index;
     n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output := n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l463_c7_2a27] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l454_c7_3583] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond;
     t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output := t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l454_c7_3583] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond;
     result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue;
     result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output := result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c7_2a27_return_output;
     VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l460_c1_87fe_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue := VAR_n_register_uxn_opcodes_phased_h_l458_c8_64e5_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l451_c7_39ed] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond;
     result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue;
     result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output := result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l451_c7_39ed] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond;
     t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output := t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l463_c1_5b59] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output;

     -- set[uxn_opcodes_phased_h_l461_c3_f77d] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l461_c3_f77d_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l461_c3_f77d_sp <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_sp;
     set_uxn_opcodes_phased_h_l461_c3_f77d_stack_index <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_stack_index;
     set_uxn_opcodes_phased_h_l461_c3_f77d_ins <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_ins;
     set_uxn_opcodes_phased_h_l461_c3_f77d_k <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_k;
     set_uxn_opcodes_phased_h_l461_c3_f77d_mul <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_mul;
     set_uxn_opcodes_phased_h_l461_c3_f77d_add <= VAR_set_uxn_opcodes_phased_h_l461_c3_f77d_add;
     -- Outputs

     -- n8_MUX[uxn_opcodes_phased_h_l457_c7_324b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_cond;
     n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output := n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l463_c1_5b59_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l457_c7_324b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l448_c2_c7e2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond;
     t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output := t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;

     -- put_stack[uxn_opcodes_phased_h_l464_c3_4b11] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l464_c3_4b11_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l464_c3_4b11_sp <= VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_sp;
     put_stack_uxn_opcodes_phased_h_l464_c3_4b11_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_stack_index;
     put_stack_uxn_opcodes_phased_h_l464_c3_4b11_offset <= VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_offset;
     put_stack_uxn_opcodes_phased_h_l464_c3_4b11_value <= VAR_put_stack_uxn_opcodes_phased_h_l464_c3_4b11_value;
     -- Outputs

     -- result_MUX[uxn_opcodes_phased_h_l448_c2_c7e2] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond;
     result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue;
     result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output := result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l454_c7_3583] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_cond;
     n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output := n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l454_c7_3583_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l451_c7_39ed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_cond;
     n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output := n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l451_c7_39ed_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l448_c2_c7e2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_cond;
     n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output := n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l448_c2_c7e2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
