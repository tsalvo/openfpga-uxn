-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity equ_0CLK_57104a4d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_57104a4d;
architecture arch of equ_0CLK_57104a4d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1229_c6_beb4]
signal BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1229_c2_b4b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1234_c11_82e7]
signal BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal n8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal t8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1234_c7_1a38]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1237_c11_c679]
signal BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1237_c7_8241]
signal n8_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1237_c7_8241]
signal t8_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1237_c7_8241]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1237_c7_8241]
signal result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1237_c7_8241]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1237_c7_8241]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1237_c7_8241]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1237_c7_8241]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1241_c11_0f1b]
signal BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1241_c7_b1e9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1244_c11_d20f]
signal BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal n8_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1244_c7_40d1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1247_c30_31fa]
signal sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1250_c21_f1f7]
signal BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1250_c21_90e8]
signal MUX_uxn_opcodes_h_l1250_c21_90e8_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1250_c21_90e8_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1250_c21_90e8_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1250_c21_90e8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1252_c11_faf0]
signal BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1252_c7_4067]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1252_c7_4067]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1252_c7_4067]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4
BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_left,
BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_right,
BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output);

-- n8_MUX_uxn_opcodes_h_l1229_c2_b4b6
n8_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- t8_MUX_uxn_opcodes_h_l1229_c2_b4b6
t8_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6
result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6
result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6
result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6
result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_left,
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_right,
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output);

-- n8_MUX_uxn_opcodes_h_l1234_c7_1a38
n8_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- t8_MUX_uxn_opcodes_h_l1234_c7_1a38
t8_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679
BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_left,
BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_right,
BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output);

-- n8_MUX_uxn_opcodes_h_l1237_c7_8241
n8_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
n8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
n8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- t8_MUX_uxn_opcodes_h_l1237_c7_8241
t8_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
t8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
t8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241
result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241
result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241
result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241
result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241
result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_left,
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_right,
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output);

-- n8_MUX_uxn_opcodes_h_l1241_c7_b1e9
n8_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f
BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_left,
BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_right,
BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output);

-- n8_MUX_uxn_opcodes_h_l1244_c7_40d1
n8_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1
result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1
result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1
result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1
result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa
sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_ins,
sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_x,
sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_y,
sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7
BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_left,
BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_right,
BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output);

-- MUX_uxn_opcodes_h_l1250_c21_90e8
MUX_uxn_opcodes_h_l1250_c21_90e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1250_c21_90e8_cond,
MUX_uxn_opcodes_h_l1250_c21_90e8_iftrue,
MUX_uxn_opcodes_h_l1250_c21_90e8_iffalse,
MUX_uxn_opcodes_h_l1250_c21_90e8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0
BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_left,
BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_right,
BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067
result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067
result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067
result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output,
 n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output,
 n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output,
 n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output,
 n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output,
 n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output,
 sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output,
 MUX_uxn_opcodes_h_l1250_c21_90e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1231_c3_999e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1235_c3_7fc3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1239_c3_6532 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1242_c3_0436 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1249_c3_2262 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1244_c7_40d1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1258_l1225_DUPLICATE_bcd3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_right := to_unsigned(5, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1235_c3_7fc3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1235_c3_7fc3;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1249_c3_2262 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1249_c3_2262;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1242_c3_0436 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1242_c3_0436;
     VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1231_c3_999e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1231_c3_999e;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1239_c3_6532 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1239_c3_6532;
     VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_iffalse := resize(to_unsigned(0, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1244_c11_d20f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1241_c11_0f1b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1237_c11_c679] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_left;
     BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output := BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1247_c30_31fa] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_ins;
     sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_x;
     sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output := sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1234_c11_82e7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1252_c11_faf0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1229_c6_beb4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1244_c7_40d1_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1250_c21_f1f7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1229_c6_beb4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_82e7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c11_c679_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_0f1b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1244_c11_d20f_return_output;
     VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1250_c21_f1f7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c11_faf0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_8c02_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1252_l1244_l1241_l1237_l1234_DUPLICATE_292e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_25d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1252_l1241_l1237_l1234_l1229_DUPLICATE_c377_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1244_l1241_l1237_l1234_l1229_DUPLICATE_d442_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1247_c30_31fa_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1252_c7_4067] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output;

     -- MUX[uxn_opcodes_h_l1250_c21_90e8] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1250_c21_90e8_cond <= VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_cond;
     MUX_uxn_opcodes_h_l1250_c21_90e8_iftrue <= VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_iftrue;
     MUX_uxn_opcodes_h_l1250_c21_90e8_iffalse <= VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_return_output := MUX_uxn_opcodes_h_l1250_c21_90e8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     t8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     t8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1252_c7_4067] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1252_c7_4067] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue := VAR_MUX_uxn_opcodes_h_l1250_c21_90e8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1252_c7_4067_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1252_c7_4067_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1252_c7_4067_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1244_c7_40d1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1244_c7_40d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     -- n8_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     n8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     n8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1241_c7_b1e9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_b1e9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- n8_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1237_c7_8241] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1237_c7_8241_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- n8_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1234_c7_1a38] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output := result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_1a38_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1229_c2_b4b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1258_l1225_DUPLICATE_bcd3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1258_l1225_DUPLICATE_bcd3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1229_c2_b4b6_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1258_l1225_DUPLICATE_bcd3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1258_l1225_DUPLICATE_bcd3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
