-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ovr_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_6d7675a8;
architecture arch of ovr_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l288_c6_65b8]
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_aae7]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l288_c2_71bc]
signal t8_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l288_c2_71bc]
signal n8_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l288_c2_71bc]
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_71bc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_71bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_71bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_71bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_71bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l289_c3_46a8[uxn_opcodes_h_l289_c3_46a8]
signal printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l293_c11_2101]
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal t8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal n8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_a4bd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l296_c11_80c0]
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l296_c7_947e]
signal t8_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l296_c7_947e]
signal n8_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l296_c7_947e]
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_947e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_947e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_947e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_947e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_947e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l299_c11_e588]
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l299_c7_777c]
signal n8_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l299_c7_777c]
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_777c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_777c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_777c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_777c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_777c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l302_c30_036c]
signal sp_relative_shift_uxn_opcodes_h_l302_c30_036c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_036c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_036c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l307_c11_0764]
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l307_c7_ede2]
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_ede2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_ede2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_ede2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_ede2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l312_c11_36a0]
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_b0e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l312_c7_b0e3]
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_b0e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_b0e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l316_c11_c915]
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_34fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_34fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8
BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_left,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_right,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output);

-- t8_MUX_uxn_opcodes_h_l288_c2_71bc
t8_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
t8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
t8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- n8_MUX_uxn_opcodes_h_l288_c2_71bc
n8_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
n8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
n8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc
result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

-- printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8
printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8 : entity work.printf_uxn_opcodes_h_l289_c3_46a8_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101
BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_left,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_right,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output);

-- t8_MUX_uxn_opcodes_h_l293_c7_a4bd
t8_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- n8_MUX_uxn_opcodes_h_l293_c7_a4bd
n8_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd
result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0
BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_left,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_right,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output);

-- t8_MUX_uxn_opcodes_h_l296_c7_947e
t8_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l296_c7_947e_cond,
t8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
t8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- n8_MUX_uxn_opcodes_h_l296_c7_947e
n8_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l296_c7_947e_cond,
n8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
n8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e
result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_cond,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588
BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_left,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_right,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output);

-- n8_MUX_uxn_opcodes_h_l299_c7_777c
n8_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l299_c7_777c_cond,
n8_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
n8_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c
result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_cond,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l302_c30_036c
sp_relative_shift_uxn_opcodes_h_l302_c30_036c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l302_c30_036c_ins,
sp_relative_shift_uxn_opcodes_h_l302_c30_036c_x,
sp_relative_shift_uxn_opcodes_h_l302_c30_036c_y,
sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_left,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_right,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2
result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_cond,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0
BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_left,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_right,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3
result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915
BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_left,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_right,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output,
 t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output,
 t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output,
 t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output,
 n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output,
 sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_dd35 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_76c4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_0856 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_815e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_df3b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_a692_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l321_l284_DUPLICATE_f6af_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_815e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_815e;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_0856 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_0856;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_76c4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_76c4;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_df3b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_df3b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_dd35 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_dd35;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l302_c30_036c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l302_c30_036c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_ins;
     sp_relative_shift_uxn_opcodes_h_l302_c30_036c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_x;
     sp_relative_shift_uxn_opcodes_h_l302_c30_036c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output := sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l312_c11_36a0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_left;
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output := BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l307_c11_0764] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_left;
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output := BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_a692 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_a692_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l299_c11_e588] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_left;
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output := BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l316_c11_c915] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_left;
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output := BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l293_c11_2101] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_left;
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output := BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l288_c6_65b8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_left;
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output := BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l296_c11_80c0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_left;
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output := BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9_return_output := result.u8_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_65b8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_2101_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_80c0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_e588_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0764_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_36a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_c915_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l288_l299_l293_l296_DUPLICATE_9c66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l293_l307_l316_l299_l312_l296_DUPLICATE_2e8d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l288_l293_l307_l296_DUPLICATE_d0f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l293_l288_l307_l316_l312_l296_DUPLICATE_3100_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_a692_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l312_l296_DUPLICATE_a692_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l288_l293_l312_l296_DUPLICATE_70c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_036c_return_output;
     -- n8_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     n8_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     n8_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output := n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- t8_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     t8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     t8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output := t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_34fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_ede2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_b0e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_34fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_aae7] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l312_c7_b0e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_aae7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_34fc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_34fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_t8_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_b0e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;

     -- n8_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     n8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     n8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output := n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_b0e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l307_c7_ede2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output := result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_ede2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;

     -- t8_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- printf_uxn_opcodes_h_l289_c3_46a8[uxn_opcodes_h_l289_c3_46a8] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l289_c3_46a8_uxn_opcodes_h_l289_c3_46a8_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_b0e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_t8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output := result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- t8_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     t8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     t8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_ede2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;

     -- n8_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_ede2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_n8_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_ede2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output := result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- n8_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     n8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     n8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_777c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_777c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_947e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_947e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_a4bd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_a4bd_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_71bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l321_l284_DUPLICATE_f6af LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l321_l284_DUPLICATE_f6af_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_71bc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_71bc_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l321_l284_DUPLICATE_f6af_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l321_l284_DUPLICATE_f6af_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
