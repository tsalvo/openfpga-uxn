-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 73
entity deo2_0CLK_5952a5d7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end deo2_0CLK_5952a5d7;
architecture arch of deo2_0CLK_5952a5d7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal current_deo_phase : unsigned(7 downto 0) := to_unsigned(0, 8);
signal deo_param0 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal deo_param1 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal is_second_deo : unsigned(0 downto 0) := to_unsigned(0, 1);
signal is_phase_3 : unsigned(0 downto 0) := to_unsigned(0, 1);
signal is_phase_4 : unsigned(0 downto 0) := to_unsigned(0, 1);
signal result : opcode_result_t := opcode_result_t_NULL;
signal device_out_result : device_out_result_t := device_out_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_current_deo_phase : unsigned(7 downto 0);
signal REG_COMB_deo_param0 : unsigned(7 downto 0);
signal REG_COMB_deo_param1 : unsigned(7 downto 0);
signal REG_COMB_is_second_deo : unsigned(0 downto 0);
signal REG_COMB_is_phase_3 : unsigned(0 downto 0);
signal REG_COMB_is_phase_4 : unsigned(0 downto 0);
signal REG_COMB_result : opcode_result_t;
signal REG_COMB_device_out_result : device_out_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l556_c6_ab6c]
signal BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l571_c7_002d]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- is_phase_4_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal n8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : device_out_result_t;

-- result_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : opcode_result_t;
signal result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : opcode_result_t;
signal result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : opcode_result_t;

-- is_phase_3_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(0 downto 0);

-- deo_param0_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal l8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal t8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l556_c2_3ba4]
signal is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l571_c11_3712]
signal BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- is_phase_4_MUX[uxn_opcodes_h_l571_c7_002d]
signal is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l571_c7_002d]
signal deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l571_c7_002d]
signal n8_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l571_c7_002d]
signal device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output : device_out_result_t;

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l571_c7_002d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(3 downto 0);

-- is_phase_3_MUX[uxn_opcodes_h_l571_c7_002d]
signal is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- deo_param0_MUX[uxn_opcodes_h_l571_c7_002d]
signal deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l571_c7_002d]
signal l8_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l571_c7_002d]
signal t8_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l571_c7_002d]
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l571_c7_002d]
signal is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l574_c11_eff5]
signal BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l578_c1_992c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output : unsigned(0 downto 0);

-- is_phase_4_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal n8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : device_out_result_t;

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(3 downto 0);

-- is_phase_3_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- deo_param0_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal l8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal t8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l574_c7_ddc0]
signal is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l579_c17_a4ce]
signal BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l579_c17_bbc8]
signal MUX_uxn_opcodes_h_l579_c17_bbc8_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l579_c17_bbc8_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l579_c17_bbc8_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l579_c17_bbc8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l580_c17_4d02]
signal BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l580_c17_2569]
signal MUX_uxn_opcodes_h_l580_c17_2569_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l580_c17_2569_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l580_c17_2569_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l580_c17_2569_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l581_c8_1c95]
signal MUX_uxn_opcodes_h_l581_c8_1c95_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l581_c8_1c95_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l581_c8_1c95_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l581_c8_1c95_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l582_c8_ec47]
signal MUX_uxn_opcodes_h_l582_c8_ec47_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l582_c8_ec47_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l582_c8_ec47_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l582_c8_ec47_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l583_c32_2d11]
signal BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output : unsigned(8 downto 0);

-- MUX[uxn_opcodes_h_l583_c16_ad6c]
signal MUX_uxn_opcodes_h_l583_c16_ad6c_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l583_c16_ad6c_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l583_c16_ad6c_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l583_c16_ad6c_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l584_c16_13c6]
signal MUX_uxn_opcodes_h_l584_c16_13c6_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l584_c16_13c6_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l584_c16_13c6_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l584_c16_13c6_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l585_c43_f403]
signal sp_relative_shift_uxn_opcodes_h_l585_c43_f403_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l585_c43_f403_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l585_c43_f403_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output : signed(3 downto 0);

-- MUX[uxn_opcodes_h_l585_c30_5996]
signal MUX_uxn_opcodes_h_l585_c30_5996_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l585_c30_5996_iftrue : signed(3 downto 0);
signal MUX_uxn_opcodes_h_l585_c30_5996_iffalse : signed(3 downto 0);
signal MUX_uxn_opcodes_h_l585_c30_5996_return_output : signed(3 downto 0);

-- device_out[uxn_opcodes_h_l586_c23_701a]
signal device_out_uxn_opcodes_h_l586_c23_701a_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_out_uxn_opcodes_h_l586_c23_701a_device_address : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l586_c23_701a_value : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l586_c23_701a_phase : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l586_c23_701a_previous_device_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l586_c23_701a_previous_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l586_c23_701a_return_output : device_out_result_t;

-- BIN_OP_AND[uxn_opcodes_h_l593_c24_9213]
signal BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_left : unsigned(0 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_right : unsigned(0 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output : unsigned(0 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l594_c3_b017]
signal current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l594_c3_b017]
signal is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l598_c4_6ab7]
signal BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4770( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.is_ram_write := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_opc_done := ref_toks_8;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a989( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_device_ram_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u16_value := ref_toks_5;
      base.device_ram_address := ref_toks_6;
      base.vram_write_layer := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c
BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_left,
BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_right,
BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4
is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4
deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- n8_MUX_uxn_opcodes_h_l556_c2_3ba4
n8_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4
device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- result_MUX_uxn_opcodes_h_l556_c2_3ba4
result_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_opcode_result_t_opcode_result_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4
is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4
deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- l8_MUX_uxn_opcodes_h_l556_c2_3ba4
l8_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- t8_MUX_uxn_opcodes_h_l556_c2_3ba4
t8_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4
current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4
is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_cond,
is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712
BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_left,
BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_right,
BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d
is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_cond,
is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l571_c7_002d
deo_param1_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_cond,
deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- n8_MUX_uxn_opcodes_h_l571_c7_002d
n8_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l571_c7_002d_cond,
n8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
n8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l571_c7_002d
device_out_result_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_cond,
device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d
result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d
result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d
result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d
result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d
result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d
result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d
result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d
result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d
is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_cond,
is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l571_c7_002d
deo_param0_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_cond,
deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- l8_MUX_uxn_opcodes_h_l571_c7_002d
l8_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l571_c7_002d_cond,
l8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
l8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- t8_MUX_uxn_opcodes_h_l571_c7_002d
t8_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l571_c7_002d_cond,
t8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
t8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d
current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_cond,
current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d
is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_cond,
is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5
BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_left,
BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_right,
BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output);

-- is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0
is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0
deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- n8_MUX_uxn_opcodes_h_l574_c7_ddc0
n8_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0
device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0
result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0
result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0
result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0
result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0
result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0
result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0
result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0
result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0
is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0
deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- l8_MUX_uxn_opcodes_h_l574_c7_ddc0
l8_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- t8_MUX_uxn_opcodes_h_l574_c7_ddc0
t8_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0
current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0
is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_cond,
is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce
BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_left,
BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_right,
BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output);

-- MUX_uxn_opcodes_h_l579_c17_bbc8
MUX_uxn_opcodes_h_l579_c17_bbc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l579_c17_bbc8_cond,
MUX_uxn_opcodes_h_l579_c17_bbc8_iftrue,
MUX_uxn_opcodes_h_l579_c17_bbc8_iffalse,
MUX_uxn_opcodes_h_l579_c17_bbc8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02
BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_left,
BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_right,
BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output);

-- MUX_uxn_opcodes_h_l580_c17_2569
MUX_uxn_opcodes_h_l580_c17_2569 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l580_c17_2569_cond,
MUX_uxn_opcodes_h_l580_c17_2569_iftrue,
MUX_uxn_opcodes_h_l580_c17_2569_iffalse,
MUX_uxn_opcodes_h_l580_c17_2569_return_output);

-- MUX_uxn_opcodes_h_l581_c8_1c95
MUX_uxn_opcodes_h_l581_c8_1c95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l581_c8_1c95_cond,
MUX_uxn_opcodes_h_l581_c8_1c95_iftrue,
MUX_uxn_opcodes_h_l581_c8_1c95_iffalse,
MUX_uxn_opcodes_h_l581_c8_1c95_return_output);

-- MUX_uxn_opcodes_h_l582_c8_ec47
MUX_uxn_opcodes_h_l582_c8_ec47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l582_c8_ec47_cond,
MUX_uxn_opcodes_h_l582_c8_ec47_iftrue,
MUX_uxn_opcodes_h_l582_c8_ec47_iffalse,
MUX_uxn_opcodes_h_l582_c8_ec47_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11
BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_left,
BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_right,
BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output);

-- MUX_uxn_opcodes_h_l583_c16_ad6c
MUX_uxn_opcodes_h_l583_c16_ad6c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l583_c16_ad6c_cond,
MUX_uxn_opcodes_h_l583_c16_ad6c_iftrue,
MUX_uxn_opcodes_h_l583_c16_ad6c_iffalse,
MUX_uxn_opcodes_h_l583_c16_ad6c_return_output);

-- MUX_uxn_opcodes_h_l584_c16_13c6
MUX_uxn_opcodes_h_l584_c16_13c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l584_c16_13c6_cond,
MUX_uxn_opcodes_h_l584_c16_13c6_iftrue,
MUX_uxn_opcodes_h_l584_c16_13c6_iffalse,
MUX_uxn_opcodes_h_l584_c16_13c6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l585_c43_f403
sp_relative_shift_uxn_opcodes_h_l585_c43_f403 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l585_c43_f403_ins,
sp_relative_shift_uxn_opcodes_h_l585_c43_f403_x,
sp_relative_shift_uxn_opcodes_h_l585_c43_f403_y,
sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output);

-- MUX_uxn_opcodes_h_l585_c30_5996
MUX_uxn_opcodes_h_l585_c30_5996 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l585_c30_5996_cond,
MUX_uxn_opcodes_h_l585_c30_5996_iftrue,
MUX_uxn_opcodes_h_l585_c30_5996_iffalse,
MUX_uxn_opcodes_h_l585_c30_5996_return_output);

-- device_out_uxn_opcodes_h_l586_c23_701a
device_out_uxn_opcodes_h_l586_c23_701a : entity work.device_out_0CLK_1666823b port map (
clk,
device_out_uxn_opcodes_h_l586_c23_701a_CLOCK_ENABLE,
device_out_uxn_opcodes_h_l586_c23_701a_device_address,
device_out_uxn_opcodes_h_l586_c23_701a_value,
device_out_uxn_opcodes_h_l586_c23_701a_phase,
device_out_uxn_opcodes_h_l586_c23_701a_previous_device_ram_read,
device_out_uxn_opcodes_h_l586_c23_701a_previous_ram_read,
device_out_uxn_opcodes_h_l586_c23_701a_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l593_c24_9213
BIN_OP_AND_uxn_opcodes_h_l593_c24_9213 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_left,
BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_right,
BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017
current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_cond,
current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017
is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_cond,
is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7
BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_left,
BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_right,
BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 previous_ram_read,
 -- Registers
 t8,
 n8,
 l8,
 current_deo_phase,
 deo_param0,
 deo_param1,
 is_second_deo,
 is_phase_3,
 is_phase_4,
 result,
 device_out_result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output,
 is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output,
 MUX_uxn_opcodes_h_l579_c17_bbc8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output,
 MUX_uxn_opcodes_h_l580_c17_2569_return_output,
 MUX_uxn_opcodes_h_l581_c8_1c95_return_output,
 MUX_uxn_opcodes_h_l582_c8_ec47_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output,
 MUX_uxn_opcodes_h_l583_c16_ad6c_return_output,
 MUX_uxn_opcodes_h_l584_c16_13c6_return_output,
 sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output,
 MUX_uxn_opcodes_h_l585_c30_5996_return_output,
 device_out_uxn_opcodes_h_l586_c23_701a_return_output,
 BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : opcode_result_t;
 variable VAR_result_TRUE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_4770_uxn_opcodes_h_l556_c2_3ba4_return_output : opcode_result_t;
 variable VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : opcode_result_t;
 variable VAR_result_FALSE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_a989_uxn_opcodes_h_l556_c2_3ba4_return_output : opcode_result_t;
 variable VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : opcode_result_t;
 variable VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l569_c3_7b61 : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l561_c3_008b : signed(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l566_c3_1b73 : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l572_c3_06a7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l575_c3_1443 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l574_c7_ddc0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l580_c17_2569_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l580_c17_2569_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l580_c17_2569_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l580_c17_2569_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l581_c8_1c95_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l581_c8_1c95_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l581_c8_1c95_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l581_c8_1c95_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l582_c8_ec47_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l582_c8_ec47_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l582_c8_ec47_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l582_c8_ec47_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output : unsigned(8 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l584_c16_13c6_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l584_c16_13c6_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l584_c16_13c6_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l584_c16_13c6_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l585_c30_5996_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l585_c30_5996_iftrue : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l585_c30_5996_iffalse : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l585_c30_5996_return_output : signed(3 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_device_address : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_value : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_phase : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_previous_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output : device_out_result_t;
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l587_c32_7799_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l588_c31_1507_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l589_c26_a8ee_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l590_c29_b17b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l591_c22_d55d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l592_c21_dc67_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l595_c4_c30c : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l598_c4_10e3 : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2c69_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_22d5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2812_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_91e0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_656c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_c216_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_cebf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_768a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l593_l594_DUPLICATE_1365_return_output : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_current_deo_phase : unsigned(7 downto 0);
variable REG_VAR_deo_param0 : unsigned(7 downto 0);
variable REG_VAR_deo_param1 : unsigned(7 downto 0);
variable REG_VAR_is_second_deo : unsigned(0 downto 0);
variable REG_VAR_is_phase_3 : unsigned(0 downto 0);
variable REG_VAR_is_phase_4 : unsigned(0 downto 0);
variable REG_VAR_result : opcode_result_t;
variable REG_VAR_device_out_result : device_out_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_current_deo_phase := current_deo_phase;
  REG_VAR_deo_param0 := deo_param0;
  REG_VAR_deo_param1 := deo_param1;
  REG_VAR_is_second_deo := is_second_deo;
  REG_VAR_is_phase_3 := is_phase_3;
  REG_VAR_is_phase_4 := is_phase_4;
  REG_VAR_result := result;
  REG_VAR_device_out_result := device_out_result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_current_deo_phase_uxn_opcodes_h_l569_c3_7b61 := resize(to_unsigned(0, 1), 8);
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := VAR_current_deo_phase_uxn_opcodes_h_l569_c3_7b61;
     VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_iftrue := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l572_c3_06a7 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l572_c3_06a7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_right := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_right := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l585_c30_5996_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_MUX_uxn_opcodes_h_l580_c17_2569_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l561_c3_008b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l575_c3_1443 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l575_c3_1443;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_y := resize(to_signed(-3, 3), 4);
     VAR_current_deo_phase_uxn_opcodes_h_l595_c4_c30c := resize(to_unsigned(0, 1), 8);
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iftrue := VAR_current_deo_phase_uxn_opcodes_h_l595_c4_c30c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l566_c3_1b73 := resize(to_unsigned(1, 1), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_right := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_right := to_unsigned(1, 1);
     VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l580_c17_2569_iffalse := to_unsigned(0, 1);
     VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_left := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := current_deo_phase;
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_phase := current_deo_phase;
     VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := deo_param0;
     VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := deo_param1;
     VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := device_out_result;
     VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_ins := VAR_ins;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := is_phase_3;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := is_phase_3;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := is_phase_3;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := is_phase_4;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := is_phase_4;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := is_phase_4;
     VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_right := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_cond := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l584_c16_13c6_cond := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iffalse := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l581_c8_1c95_iffalse := l8;
     VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := l8;
     VAR_MUX_uxn_opcodes_h_l582_c8_ec47_iffalse := n8;
     VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_left := VAR_phase;
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_previous_ram_read := VAR_previous_ram_read;
     VAR_MUX_uxn_opcodes_h_l581_c8_1c95_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l582_c8_ec47_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_left := t8;
     VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := t8;
     -- BIN_OP_PLUS[uxn_opcodes_h_l598_c4_6ab7] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_left;
     BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output := BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l585_c43_f403] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l585_c43_f403_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_ins;
     sp_relative_shift_uxn_opcodes_h_l585_c43_f403_x <= VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_x;
     sp_relative_shift_uxn_opcodes_h_l585_c43_f403_y <= VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output := sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_cebf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_cebf_return_output := result.vram_write_layer;

     -- result_TRUE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_4770[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     VAR_result_TRUE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_4770_uxn_opcodes_h_l556_c2_3ba4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4770(
     result,
     to_unsigned(0, 1),
     VAR_result_sp_relative_shift_uxn_opcodes_h_l561_c3_008b,
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l566_c3_1b73,
     to_unsigned(0, 1));

     -- BIN_OP_EQ[uxn_opcodes_h_l580_c17_4d02] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_left;
     BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output := BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l579_c17_a4ce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_left;
     BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output := BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_656c LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_656c_return_output := result.u16_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2812 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2812_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2c69 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2c69_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_768a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_768a_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l574_c11_eff5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_left;
     BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output := BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l583_c32_2d11] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_left;
     BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output := BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_22d5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_22d5_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_91e0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_91e0_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l556_c6_ab6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_c216 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_c216_return_output := result.device_ram_address;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l574_c7_ddc0_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l571_c11_3712] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_left;
     BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output := BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c6_ab6c_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l571_c11_3712_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l574_c11_eff5_return_output;
     VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l579_c17_a4ce_return_output;
     VAR_MUX_uxn_opcodes_h_l580_c17_2569_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l580_c17_4d02_return_output;
     VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_iftrue := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l583_c32_2d11_return_output, 8);
     VAR_current_deo_phase_uxn_opcodes_h_l598_c4_10e3 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l598_c4_6ab7_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_768a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_768a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_656c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_656c_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2c69_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2c69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_91e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_91e0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_22d5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_22d5_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_cebf_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_cebf_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_c216_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_c216_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2812_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l571_l574_DUPLICATE_2812_return_output;
     VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue := VAR_result_TRUE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_4770_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_MUX_uxn_opcodes_h_l585_c30_5996_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l585_c43_f403_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iffalse := VAR_current_deo_phase_uxn_opcodes_h_l598_c4_10e3;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- t8_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- MUX[uxn_opcodes_h_l580_c17_2569] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l580_c17_2569_cond <= VAR_MUX_uxn_opcodes_h_l580_c17_2569_cond;
     MUX_uxn_opcodes_h_l580_c17_2569_iftrue <= VAR_MUX_uxn_opcodes_h_l580_c17_2569_iftrue;
     MUX_uxn_opcodes_h_l580_c17_2569_iffalse <= VAR_MUX_uxn_opcodes_h_l580_c17_2569_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l580_c17_2569_return_output := MUX_uxn_opcodes_h_l580_c17_2569_return_output;

     -- MUX[uxn_opcodes_h_l583_c16_ad6c] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l583_c16_ad6c_cond <= VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_cond;
     MUX_uxn_opcodes_h_l583_c16_ad6c_iftrue <= VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_iftrue;
     MUX_uxn_opcodes_h_l583_c16_ad6c_iffalse <= VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_return_output := MUX_uxn_opcodes_h_l583_c16_ad6c_return_output;

     -- MUX[uxn_opcodes_h_l579_c17_bbc8] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l579_c17_bbc8_cond <= VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_cond;
     MUX_uxn_opcodes_h_l579_c17_bbc8_iftrue <= VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_iftrue;
     MUX_uxn_opcodes_h_l579_c17_bbc8_iffalse <= VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_return_output := MUX_uxn_opcodes_h_l579_c17_bbc8_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_MUX_uxn_opcodes_h_l581_c8_1c95_cond := VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_return_output;
     VAR_MUX_uxn_opcodes_h_l585_c30_5996_cond := VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l579_c17_bbc8_return_output;
     VAR_MUX_uxn_opcodes_h_l582_c8_ec47_cond := VAR_MUX_uxn_opcodes_h_l580_c17_2569_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l580_c17_2569_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_return_output;
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_device_address := VAR_MUX_uxn_opcodes_h_l583_c16_ad6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     -- deo_param0_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- is_phase_4_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- t8_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     t8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     t8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output := t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- MUX[uxn_opcodes_h_l585_c30_5996] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l585_c30_5996_cond <= VAR_MUX_uxn_opcodes_h_l585_c30_5996_cond;
     MUX_uxn_opcodes_h_l585_c30_5996_iftrue <= VAR_MUX_uxn_opcodes_h_l585_c30_5996_iftrue;
     MUX_uxn_opcodes_h_l585_c30_5996_iffalse <= VAR_MUX_uxn_opcodes_h_l585_c30_5996_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l585_c30_5996_return_output := MUX_uxn_opcodes_h_l585_c30_5996_return_output;

     -- MUX[uxn_opcodes_h_l582_c8_ec47] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l582_c8_ec47_cond <= VAR_MUX_uxn_opcodes_h_l582_c8_ec47_cond;
     MUX_uxn_opcodes_h_l582_c8_ec47_iftrue <= VAR_MUX_uxn_opcodes_h_l582_c8_ec47_iftrue;
     MUX_uxn_opcodes_h_l582_c8_ec47_iffalse <= VAR_MUX_uxn_opcodes_h_l582_c8_ec47_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l582_c8_ec47_return_output := MUX_uxn_opcodes_h_l582_c8_ec47_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- is_phase_3_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- MUX[uxn_opcodes_h_l581_c8_1c95] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l581_c8_1c95_cond <= VAR_MUX_uxn_opcodes_h_l581_c8_1c95_cond;
     MUX_uxn_opcodes_h_l581_c8_1c95_iftrue <= VAR_MUX_uxn_opcodes_h_l581_c8_1c95_iftrue;
     MUX_uxn_opcodes_h_l581_c8_1c95_iffalse <= VAR_MUX_uxn_opcodes_h_l581_c8_1c95_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l581_c8_1c95_return_output := MUX_uxn_opcodes_h_l581_c8_1c95_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_MUX_uxn_opcodes_h_l584_c16_13c6_iffalse := VAR_MUX_uxn_opcodes_h_l581_c8_1c95_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l581_c8_1c95_return_output;
     VAR_MUX_uxn_opcodes_h_l584_c16_13c6_iftrue := VAR_MUX_uxn_opcodes_h_l582_c8_ec47_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l582_c8_ec47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l585_c30_5996_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_is_phase_3_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_is_phase_4_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- is_phase_3_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output := is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- MUX[uxn_opcodes_h_l584_c16_13c6] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l584_c16_13c6_cond <= VAR_MUX_uxn_opcodes_h_l584_c16_13c6_cond;
     MUX_uxn_opcodes_h_l584_c16_13c6_iftrue <= VAR_MUX_uxn_opcodes_h_l584_c16_13c6_iftrue;
     MUX_uxn_opcodes_h_l584_c16_13c6_iffalse <= VAR_MUX_uxn_opcodes_h_l584_c16_13c6_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l584_c16_13c6_return_output := MUX_uxn_opcodes_h_l584_c16_13c6_return_output;

     -- t8_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- is_phase_4_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output := is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output := deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- n8_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l578_c1_992c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output;

     -- l8_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- Submodule level 4
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l578_c1_992c_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_MUX_uxn_opcodes_h_l584_c16_13c6_return_output;
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_value := VAR_MUX_uxn_opcodes_h_l584_c16_13c6_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_is_phase_3_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_is_phase_4_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_l8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     -- deo_param1_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- is_phase_3_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- n8_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     n8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     n8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output := n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- device_out[uxn_opcodes_h_l586_c23_701a] LATENCY=0
     -- Clock enable
     device_out_uxn_opcodes_h_l586_c23_701a_CLOCK_ENABLE <= VAR_device_out_uxn_opcodes_h_l586_c23_701a_CLOCK_ENABLE;
     -- Inputs
     device_out_uxn_opcodes_h_l586_c23_701a_device_address <= VAR_device_out_uxn_opcodes_h_l586_c23_701a_device_address;
     device_out_uxn_opcodes_h_l586_c23_701a_value <= VAR_device_out_uxn_opcodes_h_l586_c23_701a_value;
     device_out_uxn_opcodes_h_l586_c23_701a_phase <= VAR_device_out_uxn_opcodes_h_l586_c23_701a_phase;
     device_out_uxn_opcodes_h_l586_c23_701a_previous_device_ram_read <= VAR_device_out_uxn_opcodes_h_l586_c23_701a_previous_device_ram_read;
     device_out_uxn_opcodes_h_l586_c23_701a_previous_ram_read <= VAR_device_out_uxn_opcodes_h_l586_c23_701a_previous_ram_read;
     -- Outputs
     VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output := device_out_uxn_opcodes_h_l586_c23_701a_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- l8_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     l8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     l8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output := l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- is_phase_4_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- Submodule level 5
     REG_VAR_deo_param0 := VAR_deo_param0_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output;
     REG_VAR_is_phase_3 := VAR_is_phase_3_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     REG_VAR_is_phase_4 := VAR_is_phase_4_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_l8_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     -- deo_param1_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output := deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- l8_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d[uxn_opcodes_h_l589_c26_a8ee] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l589_c26_a8ee_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.is_vram_write;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l587_c32_7799] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l587_c32_7799_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.is_device_ram_write;

     -- n8_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d[uxn_opcodes_h_l592_c21_dc67] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l592_c21_dc67_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.u8_value;

     -- CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d[uxn_opcodes_h_l591_c22_d55d] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l591_c22_d55d_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.u16_addr;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l593_l594_DUPLICATE_1365 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l593_l594_DUPLICATE_1365_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.is_deo_done;

     -- CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d[uxn_opcodes_h_l590_c29_b17b] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l590_c29_b17b_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.vram_write_layer;

     -- CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d[uxn_opcodes_h_l588_c31_1507] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l588_c31_1507_return_output := VAR_device_out_uxn_opcodes_h_l586_c23_701a_return_output.device_ram_address;

     -- Submodule level 6
     VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l591_c22_d55d_return_output;
     VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_left := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l593_l594_DUPLICATE_1365_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_cond := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l593_l594_DUPLICATE_1365_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_cond := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l593_l594_DUPLICATE_1365_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l587_c32_7799_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l589_c26_a8ee_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l590_c29_b17b_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l588_c31_1507_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l592_c21_dc67_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     -- is_second_deo_MUX[uxn_opcodes_h_l594_c3_b017] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_cond;
     is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output := is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l593_c24_9213] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_left;
     BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output := BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output := device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l594_c3_b017] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output := current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_BIN_OP_AND_uxn_opcodes_h_l593_c24_9213_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l594_c3_b017_return_output;
     REG_VAR_deo_param1 := VAR_deo_param1_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l594_c3_b017_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l574_c7_ddc0] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output := current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- Submodule level 8
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     REG_VAR_device_out_result := VAR_device_out_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l574_c7_ddc0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output := is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l571_c7_002d] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output := current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output;

     -- Submodule level 9
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c7_002d_return_output;
     -- current_deo_phase_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- result_FALSE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_a989[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     VAR_result_FALSE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_a989_uxn_opcodes_h_l556_c2_3ba4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a989(
     result,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l571_c7_002d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l571_c7_002d_return_output);

     -- is_second_deo_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- Submodule level 10
     REG_VAR_current_deo_phase := VAR_current_deo_phase_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     REG_VAR_is_second_deo := VAR_is_second_deo_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse := VAR_result_FALSE_INPUT_MUX_CONST_REF_RD_opcode_result_t_opcode_result_t_a989_uxn_opcodes_h_l556_c2_3ba4_return_output;
     -- result_MUX[uxn_opcodes_h_l556_c2_3ba4] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond <= VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_cond;
     result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue <= VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iftrue;
     result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse <= VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output := result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;

     -- Submodule level 11
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_h_l556_c2_3ba4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_current_deo_phase <= REG_VAR_current_deo_phase;
REG_COMB_deo_param0 <= REG_VAR_deo_param0;
REG_COMB_deo_param1 <= REG_VAR_deo_param1;
REG_COMB_is_second_deo <= REG_VAR_is_second_deo;
REG_COMB_is_phase_3 <= REG_VAR_is_phase_3;
REG_COMB_is_phase_4 <= REG_VAR_is_phase_4;
REG_COMB_result <= REG_VAR_result;
REG_COMB_device_out_result <= REG_VAR_device_out_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     current_deo_phase <= REG_COMB_current_deo_phase;
     deo_param0 <= REG_COMB_deo_param0;
     deo_param1 <= REG_COMB_deo_param1;
     is_second_deo <= REG_COMB_is_second_deo;
     is_phase_3 <= REG_COMB_is_phase_3;
     is_phase_4 <= REG_COMB_is_phase_4;
     result <= REG_COMB_result;
     device_out_result <= REG_COMB_device_out_result;
 end if;
 end if;
end process;

end arch;
