-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity opc_equ_phased_0CLK_2ca51e56 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_equ_phased_0CLK_2ca51e56;
architecture arch of opc_equ_phased_0CLK_2ca51e56 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l418_c6_14f4]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l418_c1_fbd6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l421_c7_35d4]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l418_c2_bf8d]
signal t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l418_c2_bf8d]
signal n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l418_c2_bf8d]
signal result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l419_c12_5a73]
signal set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l421_c11_f99e]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l421_c1_c695]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l424_c7_9843]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l421_c7_35d4]
signal t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l421_c7_35d4]
signal n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l421_c7_35d4]
signal result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l422_c8_86b4]
signal t_register_uxn_opcodes_phased_h_l422_c8_86b4_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l424_c11_b021]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l424_c1_a2e6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l427_c7_2c67]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l424_c7_9843]
signal t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l424_c7_9843]
signal n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l424_c7_9843]
signal result_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l425_c8_a381]
signal n_register_uxn_opcodes_phased_h_l425_c8_a381_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l427_c11_a500]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l427_c1_7c36]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l430_c7_7b31]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l427_c7_2c67]
signal n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l427_c7_2c67]
signal result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l428_c8_12ed]
signal n_register_uxn_opcodes_phased_h_l428_c8_12ed_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l430_c11_8f6f]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l430_c1_b560]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l433_c7_9110]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l430_c7_7b31]
signal result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l431_c3_6a1b]
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l431_c3_6a1b_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l433_c11_8cbb]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l433_c1_78d8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l433_c7_9110]
signal result_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l434_c33_f683]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_phased_h_l434_c33_72ed]
signal MUX_uxn_opcodes_phased_h_l434_c33_72ed_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_phased_h_l434_c33_72ed_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_phased_h_l434_c33_72ed_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_phased_h_l434_c3_74d3]
signal put_stack_uxn_opcodes_phased_h_l434_c3_74d3_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l434_c3_74d3_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l434_c3_74d3_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l434_c3_74d3_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l434_c3_74d3_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l436_c11_970c]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l436_c7_00fd]
signal result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4
BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d
t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond,
t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue,
t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse,
t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d
n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond,
n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue,
n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse,
n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output);

-- result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d
result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond,
result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue,
result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse,
result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_sp,
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_k,
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_mul,
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_add,
set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e
BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4
t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond,
t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue,
t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse,
t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4
n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond,
n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue,
n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse,
n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output);

-- result_MUX_uxn_opcodes_phased_h_l421_c7_35d4
result_MUX_uxn_opcodes_phased_h_l421_c7_35d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond,
result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue,
result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse,
result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output);

-- t_register_uxn_opcodes_phased_h_l422_c8_86b4
t_register_uxn_opcodes_phased_h_l422_c8_86b4 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l422_c8_86b4_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_index,
t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_ptr,
t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021
BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l424_c7_9843
t8_MUX_uxn_opcodes_phased_h_l424_c7_9843 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond,
t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue,
t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse,
t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l424_c7_9843
n8_MUX_uxn_opcodes_phased_h_l424_c7_9843 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond,
n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue,
n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse,
n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output);

-- result_MUX_uxn_opcodes_phased_h_l424_c7_9843
result_MUX_uxn_opcodes_phased_h_l424_c7_9843 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond,
result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue,
result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse,
result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output);

-- n_register_uxn_opcodes_phased_h_l425_c8_a381
n_register_uxn_opcodes_phased_h_l425_c8_a381 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l425_c8_a381_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_index,
n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_ptr,
n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500
BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67
n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond,
n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue,
n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse,
n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output);

-- result_MUX_uxn_opcodes_phased_h_l427_c7_2c67
result_MUX_uxn_opcodes_phased_h_l427_c7_2c67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond,
result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue,
result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse,
result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output);

-- n_register_uxn_opcodes_phased_h_l428_c8_12ed
n_register_uxn_opcodes_phased_h_l428_c8_12ed : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l428_c8_12ed_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_index,
n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_ptr,
n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f
BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output);

-- result_MUX_uxn_opcodes_phased_h_l430_c7_7b31
result_MUX_uxn_opcodes_phased_h_l430_c7_7b31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond,
result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue,
result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse,
result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output);

-- set_uxn_opcodes_phased_h_l431_c3_6a1b
set_uxn_opcodes_phased_h_l431_c3_6a1b : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l431_c3_6a1b_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l431_c3_6a1b_sp,
set_uxn_opcodes_phased_h_l431_c3_6a1b_stack_index,
set_uxn_opcodes_phased_h_l431_c3_6a1b_ins,
set_uxn_opcodes_phased_h_l431_c3_6a1b_k,
set_uxn_opcodes_phased_h_l431_c3_6a1b_mul,
set_uxn_opcodes_phased_h_l431_c3_6a1b_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb
BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output);

-- result_MUX_uxn_opcodes_phased_h_l433_c7_9110
result_MUX_uxn_opcodes_phased_h_l433_c7_9110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond,
result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue,
result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse,
result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683
BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output);

-- MUX_uxn_opcodes_phased_h_l434_c33_72ed
MUX_uxn_opcodes_phased_h_l434_c33_72ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_phased_h_l434_c33_72ed_cond,
MUX_uxn_opcodes_phased_h_l434_c33_72ed_iftrue,
MUX_uxn_opcodes_phased_h_l434_c33_72ed_iffalse,
MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output);

-- put_stack_uxn_opcodes_phased_h_l434_c3_74d3
put_stack_uxn_opcodes_phased_h_l434_c3_74d3 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l434_c3_74d3_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l434_c3_74d3_sp,
put_stack_uxn_opcodes_phased_h_l434_c3_74d3_stack_index,
put_stack_uxn_opcodes_phased_h_l434_c3_74d3_offset,
put_stack_uxn_opcodes_phased_h_l434_c3_74d3_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c
BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l436_c7_00fd
result_MUX_uxn_opcodes_phased_h_l436_c7_00fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_cond,
result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iftrue,
result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iffalse,
result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output,
 t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output,
 n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output,
 result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output,
 set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output,
 t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output,
 n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output,
 result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output,
 t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output,
 t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output,
 n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output,
 result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output,
 n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output,
 n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output,
 result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output,
 n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output,
 result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output,
 result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output,
 MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output,
 result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_value : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_add := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_right := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_right := to_unsigned(6, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue := to_unsigned(0, 1);
     VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_offset := resize(to_unsigned(0, 1), 8);
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_add := resize(to_signed(-1, 2), 8);
     VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_k := VAR_k;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_index := VAR_stack_index;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_right := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l430_c11_8f6f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l436_c11_970c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l427_c11_a500] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l433_c11_8cbb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l421_c11_f99e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l418_c6_14f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l434_c33_f683] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l424_c11_b021] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l418_c6_14f4_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l421_c11_f99e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l424_c11_b021_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l427_c11_a500_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l430_c11_8f6f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l433_c11_8cbb_return_output;
     VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l434_c33_f683_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l436_c11_970c_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l421_c7_35d4] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l418_c1_fbd6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l436_c7_00fd] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_cond;
     result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iftrue;
     result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output := result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output;

     -- MUX[uxn_opcodes_phased_h_l434_c33_72ed] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_phased_h_l434_c33_72ed_cond <= VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_cond;
     MUX_uxn_opcodes_phased_h_l434_c33_72ed_iftrue <= VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_iftrue;
     MUX_uxn_opcodes_phased_h_l434_c33_72ed_iffalse <= VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output := MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_value := VAR_MUX_uxn_opcodes_phased_h_l434_c33_72ed_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l418_c1_fbd6_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l436_c7_00fd_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l424_c7_9843] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l433_c7_9110] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond;
     result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue;
     result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output := result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l421_c1_c695] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l419_c12_5a73] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_sp;
     set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_k;
     set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_mul;
     set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output := set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l421_c1_c695_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l419_c12_5a73_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l427_c7_2c67] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l430_c7_7b31] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond;
     result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue;
     result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output := result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output;

     -- t_register[uxn_opcodes_phased_h_l422_c8_86b4] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l422_c8_86b4_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_index;
     t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output := t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l424_c1_a2e6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l424_c1_a2e6_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue := VAR_t_register_uxn_opcodes_phased_h_l422_c8_86b4_return_output;
     -- n_register[uxn_opcodes_phased_h_l425_c8_a381] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l425_c8_a381_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_index;
     n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output := n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l430_c7_7b31] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l427_c7_2c67] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond;
     result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue;
     result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output := result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l427_c1_7c36] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c7_7b31_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l427_c1_7c36_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue := VAR_n_register_uxn_opcodes_phased_h_l425_c8_a381_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l424_c7_9843] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond;
     result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue;
     result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output := result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l430_c1_b560] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l424_c7_9843] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond;
     t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output := t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l433_c7_9110] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output;

     -- n_register[uxn_opcodes_phased_h_l428_c8_12ed] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l428_c8_12ed_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_index;
     n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output := n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c7_9110_return_output;
     VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l430_c1_b560_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue := VAR_n_register_uxn_opcodes_phased_h_l428_c8_12ed_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;
     -- set[uxn_opcodes_phased_h_l431_c3_6a1b] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l431_c3_6a1b_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l431_c3_6a1b_sp <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_sp;
     set_uxn_opcodes_phased_h_l431_c3_6a1b_stack_index <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_stack_index;
     set_uxn_opcodes_phased_h_l431_c3_6a1b_ins <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_ins;
     set_uxn_opcodes_phased_h_l431_c3_6a1b_k <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_k;
     set_uxn_opcodes_phased_h_l431_c3_6a1b_mul <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_mul;
     set_uxn_opcodes_phased_h_l431_c3_6a1b_add <= VAR_set_uxn_opcodes_phased_h_l431_c3_6a1b_add;
     -- Outputs

     -- t8_MUX[uxn_opcodes_phased_h_l421_c7_35d4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond;
     t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output := t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l421_c7_35d4] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond;
     result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue;
     result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output := result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l427_c7_2c67] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_cond;
     n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output := n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l433_c1_78d8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output;

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l433_c1_78d8_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l427_c7_2c67_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l418_c2_bf8d] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond;
     result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue;
     result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output := result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l418_c2_bf8d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond;
     t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output := t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;

     -- put_stack[uxn_opcodes_phased_h_l434_c3_74d3] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l434_c3_74d3_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l434_c3_74d3_sp <= VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_sp;
     put_stack_uxn_opcodes_phased_h_l434_c3_74d3_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_stack_index;
     put_stack_uxn_opcodes_phased_h_l434_c3_74d3_offset <= VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_offset;
     put_stack_uxn_opcodes_phased_h_l434_c3_74d3_value <= VAR_put_stack_uxn_opcodes_phased_h_l434_c3_74d3_value;
     -- Outputs

     -- n8_MUX[uxn_opcodes_phased_h_l424_c7_9843] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_cond;
     n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output := n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l424_c7_9843_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l421_c7_35d4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_cond;
     n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output := n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l421_c7_35d4_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l418_c2_bf8d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_cond;
     n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output := n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l418_c2_bf8d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
