-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity ldr_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_f74745d5;
architecture arch of ldr_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1622_c6_1180]
signal BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal t8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1622_c2_99b9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1635_c11_549d]
signal BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal t8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1635_c7_fb65]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1638_c11_85fa]
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1638_c7_6601]
signal t8_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1638_c7_6601]
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1638_c7_6601]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1638_c7_6601]
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1638_c7_6601]
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1638_c7_6601]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1638_c7_6601]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1638_c7_6601]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1640_c30_af6e]
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1641_c22_e2f9]
signal BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1643_c11_01ec]
signal BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1643_c7_eaca]
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1643_c7_eaca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1643_c7_eaca]
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1643_c7_eaca]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1643_c7_eaca]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1643_c7_eaca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1646_c11_ddb9]
signal BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1646_c7_3db9]
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1646_c7_3db9]
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1646_c7_3db9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1646_c7_3db9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1646_c7_3db9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_1a75( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;
      base.is_pc_updated := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_left,
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_right,
BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output);

-- t8_MUX_uxn_opcodes_h_l1622_c2_99b9
t8_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9
tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_left,
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_right,
BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output);

-- t8_MUX_uxn_opcodes_h_l1635_c7_fb65
t8_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65
tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_left,
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_right,
BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output);

-- t8_MUX_uxn_opcodes_h_l1638_c7_6601
t8_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
t8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
t8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1638_c7_6601
tmp8_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e
sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_ins,
sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_x,
sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_y,
sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_left,
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_right,
BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_left,
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_right,
BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca
tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_cond,
tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue,
tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse,
tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_cond,
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_left,
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_right,
BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9
tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_cond,
tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue,
tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse,
tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output,
 t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output,
 t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output,
 t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output,
 sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output,
 tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output,
 tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1627_c3_b935 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1632_c3_f9fc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1636_c3_e849 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1641_c3_13d7 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1641_c27_0f03_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1644_c3_39fc : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1649_c3_01d3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1635_l1638_l1622_DUPLICATE_703f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1635_l1643_DUPLICATE_9727_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1646_l1638_l1643_DUPLICATE_b4bf_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l1618_l1654_DUPLICATE_36f7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1644_c3_39fc := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1644_c3_39fc;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1632_c3_f9fc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1632_c3_f9fc;
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1649_c3_01d3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1649_c3_01d3;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1636_c3_e849 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1636_c3_e849;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1627_c3_b935 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1627_c3_b935;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1638_c11_85fa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_left;
     BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output := BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1643_c11_01ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1635_l1643_DUPLICATE_9727 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1635_l1643_DUPLICATE_9727_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1635_c11_549d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1640_c30_af6e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_ins;
     sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_x;
     sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output := sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1641_c27_0f03] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1641_c27_0f03_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1646_c11_ddb9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1646_l1638_l1643_DUPLICATE_b4bf LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1646_l1638_l1643_DUPLICATE_b4bf_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1635_l1638_l1622_DUPLICATE_703f LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1635_l1638_l1622_DUPLICATE_703f_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1622_c6_1180] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_left;
     BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output := BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1622_c6_1180_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1635_c11_549d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c11_85fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1643_c11_01ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1646_c11_ddb9_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1641_c27_0f03_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1635_l1643_DUPLICATE_9727_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1635_l1643_DUPLICATE_9727_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1635_l1638_l1622_DUPLICATE_703f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1635_l1638_l1622_DUPLICATE_703f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1635_l1638_l1622_DUPLICATE_703f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_7b9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1635_l1646_l1638_l1643_DUPLICATE_f79d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1646_l1638_l1643_DUPLICATE_b4bf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1646_l1638_l1643_DUPLICATE_b4bf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1646_l1638_l1643_DUPLICATE_b4bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1646_l1643_l1638_l1635_l1622_DUPLICATE_2e4a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1622_c2_99b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1640_c30_af6e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1643_c7_eaca] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;

     -- t8_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     t8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     t8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1646_c7_3db9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1646_c7_3db9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1646_c7_3db9] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_cond;
     tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output := tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1641_c22_e2f9] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1646_c7_3db9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1646_c7_3db9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1641_c3_13d7 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1641_c22_e2f9_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1646_c7_3db9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1641_c3_13d7;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1643_c7_eaca] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1643_c7_eaca] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output := result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;

     -- t8_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1643_c7_eaca] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_cond;
     tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output := tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1643_c7_eaca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1643_c7_eaca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1643_c7_eaca_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- t8_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1638_c7_6601] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1638_c7_6601_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1635_c7_fb65] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_cond;
     tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output := tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1635_c7_fb65_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1622_c2_99b9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l1618_l1654_DUPLICATE_36f7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l1618_l1654_DUPLICATE_36f7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1a75(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1622_c2_99b9_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l1618_l1654_DUPLICATE_36f7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l1618_l1654_DUPLICATE_36f7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
