-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity sth_0CLK_d6c995e8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_d6c995e8;
architecture arch of sth_0CLK_d6c995e8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2597_c6_d0d0]
signal BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2597_c1_a0b2]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2597_c2_a2b8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2598_c3_b784[uxn_opcodes_h_l2598_c3_b784]
signal printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2602_c11_0125]
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2602_c7_e9fd]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2605_c11_249f]
signal BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2605_c7_f393]
signal t8_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2605_c7_f393]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2608_c32_1373]
signal BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2608_c32_819b]
signal BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2608_c32_482e]
signal MUX_uxn_opcodes_h_l2608_c32_482e_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2608_c32_482e_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2608_c32_482e_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2608_c32_482e_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2610_c11_1544]
signal BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2610_c7_3509]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2614_c11_c5c5]
signal BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2614_c7_6b9e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2614_c7_6b9e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2614_c7_6b9e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2614_c7_6b9e]
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2614_c7_6b9e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2614_c7_6b9e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2620_c11_3363]
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2620_c7_c2b4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2620_c7_c2b4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2620_c7_c2b4]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_06e4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_value := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.is_stack_index_flipped := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0
BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_left,
BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_right,
BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output);

-- t8_MUX_uxn_opcodes_h_l2597_c2_a2b8
t8_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

-- printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784
printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784 : entity work.printf_uxn_opcodes_h_l2598_c3_b784_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125
BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_left,
BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_right,
BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output);

-- t8_MUX_uxn_opcodes_h_l2602_c7_e9fd
t8_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f
BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_left,
BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_right,
BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output);

-- t8_MUX_uxn_opcodes_h_l2605_c7_f393
t8_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
t8_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
t8_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393
result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393
result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393
result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393
result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393
result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373
BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_left,
BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_right,
BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b
BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_left,
BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_right,
BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output);

-- MUX_uxn_opcodes_h_l2608_c32_482e
MUX_uxn_opcodes_h_l2608_c32_482e : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2608_c32_482e_cond,
MUX_uxn_opcodes_h_l2608_c32_482e_iftrue,
MUX_uxn_opcodes_h_l2608_c32_482e_iffalse,
MUX_uxn_opcodes_h_l2608_c32_482e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544
BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_left,
BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_right,
BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509
result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509
result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509
result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509
result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509
result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_left,
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_right,
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond,
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363
BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_left,
BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_right,
BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output,
 t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output,
 t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output,
 t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output,
 MUX_uxn_opcodes_h_l2608_c32_482e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2599_c3_b1a5 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2603_c3_6555 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2608_c32_482e_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2608_c32_482e_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2608_c32_482e_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2608_c32_482e_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2612_c3_db4f : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2617_c3_6d26 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2597_l2610_l2602_DUPLICATE_a8be_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2614_l2605_l2610_DUPLICATE_6321_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_06e4_uxn_opcodes_h_l2593_l2626_DUPLICATE_c285_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_right := to_unsigned(4, 3);
     VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_right := to_unsigned(128, 8);
     VAR_MUX_uxn_opcodes_h_l2608_c32_482e_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2617_c3_6d26 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2617_c3_6d26;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l2608_c32_482e_iffalse := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_right := to_unsigned(5, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2612_c3_db4f := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2612_c3_db4f;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2603_c3_6555 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2603_c3_6555;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2599_c3_b1a5 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2599_c3_b1a5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2602_c11_0125] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_left;
     BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output := BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2597_c6_d0d0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2605_c11_249f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2610_c11_1544] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_left;
     BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output := BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2614_c11_c5c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2608_c32_1373] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_left;
     BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output := BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2597_l2610_l2602_DUPLICATE_a8be LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2597_l2610_l2602_DUPLICATE_a8be_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2614_l2605_l2610_DUPLICATE_6321 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2614_l2605_l2610_DUPLICATE_6321_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2620_c11_3363] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_left;
     BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output := BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2608_c32_1373_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2597_c6_d0d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c11_0125_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2605_c11_249f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2610_c11_1544_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_c5c5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c11_3363_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2597_l2610_l2602_DUPLICATE_a8be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2597_l2610_l2602_DUPLICATE_a8be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2597_l2610_l2602_DUPLICATE_a8be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2620_DUPLICATE_cd6e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2614_l2597_l2610_l2602_DUPLICATE_3b7a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2614_l2605_l2602_l2597_l2620_DUPLICATE_ee09_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2610_l2605_l2602_l2597_l2620_DUPLICATE_6f30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2614_l2605_l2610_DUPLICATE_6321_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2614_l2605_l2610_DUPLICATE_6321_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2614_l2605_l2610_DUPLICATE_6321_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2614_l2610_l2605_l2602_l2597_DUPLICATE_aade_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2614_c7_6b9e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2608_c32_819b] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_left;
     BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output := BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     t8_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     t8_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2614_c7_6b9e] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output := result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2614_c7_6b9e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2620_c7_c2b4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2597_c1_a0b2] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2620_c7_c2b4] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2620_c7_c2b4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2608_c32_482e_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2608_c32_819b_return_output;
     VAR_printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2597_c1_a0b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c7_c2b4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2614_c7_6b9e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2614_c7_6b9e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;

     -- MUX[uxn_opcodes_h_l2608_c32_482e] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2608_c32_482e_cond <= VAR_MUX_uxn_opcodes_h_l2608_c32_482e_cond;
     MUX_uxn_opcodes_h_l2608_c32_482e_iftrue <= VAR_MUX_uxn_opcodes_h_l2608_c32_482e_iftrue;
     MUX_uxn_opcodes_h_l2608_c32_482e_iffalse <= VAR_MUX_uxn_opcodes_h_l2608_c32_482e_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2608_c32_482e_return_output := MUX_uxn_opcodes_h_l2608_c32_482e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2614_c7_6b9e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- printf_uxn_opcodes_h_l2598_c3_b784[uxn_opcodes_h_l2598_c3_b784] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2598_c3_b784_uxn_opcodes_h_l2598_c3_b784_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_value_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue := VAR_MUX_uxn_opcodes_h_l2608_c32_482e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_6b9e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- t8_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2610_c7_3509] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2610_c7_3509_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2605_c7_f393] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2605_c7_f393_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2602_c7_e9fd] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c7_e9fd_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2597_c2_a2b8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_06e4_uxn_opcodes_h_l2593_l2626_DUPLICATE_c285 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_06e4_uxn_opcodes_h_l2593_l2626_DUPLICATE_c285_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_06e4(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2597_c2_a2b8_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_06e4_uxn_opcodes_h_l2593_l2626_DUPLICATE_c285_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_06e4_uxn_opcodes_h_l2593_l2626_DUPLICATE_c285_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
