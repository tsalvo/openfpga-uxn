-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity jcn2_0CLK_12273847 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jcn2_0CLK_12273847;
architecture arch of jcn2_0CLK_12273847 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l693_c6_1571]
signal BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal t16_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l693_c2_5f9b]
signal n8_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l706_c11_bc23]
signal BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l706_c7_09e9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l706_c7_09e9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l706_c7_09e9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l706_c7_09e9]
signal result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l706_c7_09e9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l706_c7_09e9]
signal t16_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l706_c7_09e9]
signal n8_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l709_c11_fa25]
signal BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l709_c7_65da]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l709_c7_65da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l709_c7_65da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l709_c7_65da]
signal result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l709_c7_65da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l709_c7_65da]
signal t16_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l709_c7_65da]
signal n8_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l711_c3_aa55]
signal CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l714_c11_2104]
signal BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l714_c7_4da8]
signal result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l714_c7_4da8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l714_c7_4da8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l714_c7_4da8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l714_c7_4da8]
signal t16_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l714_c7_4da8]
signal n8_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l715_c3_4a5b]
signal BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l717_c11_70a6]
signal BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l717_c7_2b6e]
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l717_c7_2b6e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l717_c7_2b6e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l717_c7_2b6e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l717_c7_2b6e]
signal n8_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l719_c30_41e3]
signal sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l720_c26_425a]
signal BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l720_c26_1e08]
signal MUX_uxn_opcodes_h_l720_c26_1e08_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l720_c26_1e08_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l720_c26_1e08_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l720_c26_1e08_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l721_c22_dc31]
signal BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l721_c22_1d4a]
signal MUX_uxn_opcodes_h_l721_c22_1d4a_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l721_c22_1d4a_iftrue : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l721_c22_1d4a_iffalse : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l721_c22_1d4a_return_output : unsigned(15 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571
BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_left,
BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_right,
BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b
result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b
result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b
result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b
result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b
result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- t16_MUX_uxn_opcodes_h_l693_c2_5f9b
t16_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- n8_MUX_uxn_opcodes_h_l693_c2_5f9b
n8_MUX_uxn_opcodes_h_l693_c2_5f9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l693_c2_5f9b_cond,
n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue,
n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse,
n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23
BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_left,
BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_right,
BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9
result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9
result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- t16_MUX_uxn_opcodes_h_l706_c7_09e9
t16_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
t16_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
t16_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- n8_MUX_uxn_opcodes_h_l706_c7_09e9
n8_MUX_uxn_opcodes_h_l706_c7_09e9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l706_c7_09e9_cond,
n8_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue,
n8_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse,
n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25
BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_left,
BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_right,
BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da
result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_cond,
result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- t16_MUX_uxn_opcodes_h_l709_c7_65da
t16_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l709_c7_65da_cond,
t16_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
t16_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- n8_MUX_uxn_opcodes_h_l709_c7_65da
n8_MUX_uxn_opcodes_h_l709_c7_65da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l709_c7_65da_cond,
n8_MUX_uxn_opcodes_h_l709_c7_65da_iftrue,
n8_MUX_uxn_opcodes_h_l709_c7_65da_iffalse,
n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output);

-- CONST_SL_8_uxn_opcodes_h_l711_c3_aa55
CONST_SL_8_uxn_opcodes_h_l711_c3_aa55 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_x,
CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104
BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_left,
BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_right,
BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8
result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_cond,
result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8
result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8
result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8
result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output);

-- t16_MUX_uxn_opcodes_h_l714_c7_4da8
t16_MUX_uxn_opcodes_h_l714_c7_4da8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l714_c7_4da8_cond,
t16_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue,
t16_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse,
t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output);

-- n8_MUX_uxn_opcodes_h_l714_c7_4da8
n8_MUX_uxn_opcodes_h_l714_c7_4da8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l714_c7_4da8_cond,
n8_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue,
n8_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse,
n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b
BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_left,
BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_right,
BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6
BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_left,
BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_right,
BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e
result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_cond,
result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output);

-- n8_MUX_uxn_opcodes_h_l717_c7_2b6e
n8_MUX_uxn_opcodes_h_l717_c7_2b6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l717_c7_2b6e_cond,
n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue,
n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse,
n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l719_c30_41e3
sp_relative_shift_uxn_opcodes_h_l719_c30_41e3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_ins,
sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_x,
sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_y,
sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a
BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_left,
BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_right,
BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output);

-- MUX_uxn_opcodes_h_l720_c26_1e08
MUX_uxn_opcodes_h_l720_c26_1e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l720_c26_1e08_cond,
MUX_uxn_opcodes_h_l720_c26_1e08_iftrue,
MUX_uxn_opcodes_h_l720_c26_1e08_iffalse,
MUX_uxn_opcodes_h_l720_c26_1e08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31
BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_left,
BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_right,
BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output);

-- MUX_uxn_opcodes_h_l721_c22_1d4a
MUX_uxn_opcodes_h_l721_c22_1d4a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l721_c22_1d4a_cond,
MUX_uxn_opcodes_h_l721_c22_1d4a_iftrue,
MUX_uxn_opcodes_h_l721_c22_1d4a_iffalse,
MUX_uxn_opcodes_h_l721_c22_1d4a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output,
 CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output,
 t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output,
 n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output,
 BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output,
 n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output,
 sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output,
 MUX_uxn_opcodes_h_l720_c26_1e08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output,
 MUX_uxn_opcodes_h_l721_c22_1d4a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l698_c3_e278 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l703_c3_e273 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l707_c3_97ef : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l712_c3_b46c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l709_c7_65da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l720_c26_1e08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l720_c26_1e08_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l720_c26_1e08_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l720_c26_1e08_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_iftrue : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_iffalse : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l715_l710_DUPLICATE_bda1_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc_uxn_opcodes_h_l725_l688_DUPLICATE_83f0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l712_c3_b46c := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l712_c3_b46c;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l707_c3_97ef := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l707_c3_97ef;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_iftrue := resize(to_unsigned(0, 1), 16);
     VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l698_c3_e278 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l698_c3_e278;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l720_c26_1e08_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l720_c26_1e08_iffalse := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l703_c3_e273 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l703_c3_e273;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_left := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_left := t16;
     VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_iffalse := t16;
     VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l706_c11_bc23] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_left;
     BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output := BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l719_c30_41e3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_ins;
     sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_x;
     sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output := sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l709_c11_fa25] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_left;
     BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output := BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l721_c22_dc31] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_left;
     BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output := BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l717_c11_70a6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_left;
     BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output := BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l715_l710_DUPLICATE_bda1 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l715_l710_DUPLICATE_bda1_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l714_c11_2104] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_left;
     BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output := BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l693_c6_1571] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_left;
     BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output := BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l709_c7_65da_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l720_c26_425a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_left;
     BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output := BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c6_1571_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c11_bc23_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_fa25_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l714_c11_2104_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_70a6_return_output;
     VAR_MUX_uxn_opcodes_h_l720_c26_1e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c26_425a_return_output;
     VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c22_dc31_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l715_l710_DUPLICATE_bda1_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l715_l710_DUPLICATE_bda1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_e4e5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l714_l717_l706_l709_DUPLICATE_1547_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_5675_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l714_l706_l709_DUPLICATE_bf7d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l693_c2_5f9b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l709_c7_65da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l719_c30_41e3_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- MUX[uxn_opcodes_h_l720_c26_1e08] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l720_c26_1e08_cond <= VAR_MUX_uxn_opcodes_h_l720_c26_1e08_cond;
     MUX_uxn_opcodes_h_l720_c26_1e08_iftrue <= VAR_MUX_uxn_opcodes_h_l720_c26_1e08_iftrue;
     MUX_uxn_opcodes_h_l720_c26_1e08_iffalse <= VAR_MUX_uxn_opcodes_h_l720_c26_1e08_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l720_c26_1e08_return_output := MUX_uxn_opcodes_h_l720_c26_1e08_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l717_c7_2b6e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;

     -- MUX[uxn_opcodes_h_l721_c22_1d4a] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l721_c22_1d4a_cond <= VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_cond;
     MUX_uxn_opcodes_h_l721_c22_1d4a_iftrue <= VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_iftrue;
     MUX_uxn_opcodes_h_l721_c22_1d4a_iffalse <= VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_return_output := MUX_uxn_opcodes_h_l721_c22_1d4a_return_output;

     -- n8_MUX[uxn_opcodes_h_l717_c7_2b6e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l717_c7_2b6e_cond <= VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_cond;
     n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue;
     n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output := n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l715_c3_4a5b] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_left;
     BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output := BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l711_c3_aa55] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_x <= VAR_CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output := CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l717_c7_2b6e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l715_c3_4a5b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l711_c3_aa55_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue := VAR_MUX_uxn_opcodes_h_l720_c26_1e08_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue := VAR_MUX_uxn_opcodes_h_l721_c22_1d4a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l714_c7_4da8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;

     -- t16_MUX[uxn_opcodes_h_l714_c7_4da8] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l714_c7_4da8_cond <= VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_cond;
     t16_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue;
     t16_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output := t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l717_c7_2b6e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output := result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l717_c7_2b6e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;

     -- n8_MUX[uxn_opcodes_h_l714_c7_4da8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l714_c7_4da8_cond <= VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_cond;
     n8_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue;
     n8_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output := n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l714_c7_4da8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_n8_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_2b6e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_t16_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;
     -- t16_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     t16_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     t16_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output := t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l714_c7_4da8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output := result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- n8_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     n8_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     n8_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output := n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l714_c7_4da8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l714_c7_4da8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_t16_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     -- n8_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     n8_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     n8_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- t16_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     t16_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     t16_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l709_c7_65da] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_cond;
     result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output := result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l709_c7_65da_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_t16_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- t16_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- n8_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l706_c7_09e9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c7_09e9_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l693_c2_5f9b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc_uxn_opcodes_h_l725_l688_DUPLICATE_83f0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc_uxn_opcodes_h_l725_l688_DUPLICATE_83f0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c2_5f9b_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc_uxn_opcodes_h_l725_l688_DUPLICATE_83f0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6bdc_uxn_opcodes_h_l725_l688_DUPLICATE_83f0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
