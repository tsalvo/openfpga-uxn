-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sth_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_85d5529e;
architecture arch of sth_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2259_c6_2674]
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2259_c1_b977]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal t8_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2259_c2_fdff]
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2260_c3_d844[uxn_opcodes_h_l2260_c3_d844]
signal printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2264_c11_8ba0]
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2264_c7_535f]
signal t8_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2264_c7_535f]
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2267_c11_f905]
signal BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2267_c7_1128]
signal t8_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2267_c7_1128]
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2270_c30_3fda]
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2272_c11_860e]
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2272_c7_58e3]
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2279_c11_5867]
signal BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2279_c7_4a47]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2279_c7_4a47]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2279_c7_4a47]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2279_c7_4a47]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_12f7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.u8_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_left,
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_right,
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output);

-- t8_MUX_uxn_opcodes_h_l2259_c2_fdff
t8_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_cond,
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

-- printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844
printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844 : entity work.printf_uxn_opcodes_h_l2260_c3_d844_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_left,
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_right,
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output);

-- t8_MUX_uxn_opcodes_h_l2264_c7_535f
t8_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
t8_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
t8_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_left,
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_right,
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output);

-- t8_MUX_uxn_opcodes_h_l2267_c7_1128
t8_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
t8_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
t8_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_cond,
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda
sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_ins,
sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_x,
sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_y,
sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_left,
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_right,
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_left,
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_right,
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output,
 t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output,
 t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output,
 t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output,
 sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_2776 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2265_c3_5587 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2276_c3_5ecc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2274_c3_cfb3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_DUPLICATE_20ea_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2272_l2267_DUPLICATE_2f87_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_12f7_uxn_opcodes_h_l2286_l2255_DUPLICATE_90ee_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_right := to_unsigned(4, 3);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2276_c3_5ecc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2276_c3_5ecc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2265_c3_5587 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2265_c3_5587;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2274_c3_cfb3 := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2274_c3_cfb3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_2776 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_2776;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2272_c11_860e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2259_c6_2674] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_left;
     BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output := BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2279_c11_5867] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_left;
     BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output := BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2264_c11_8ba0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2267_c11_f905] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_left;
     BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output := BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2270_c30_3fda] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_ins;
     sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_x;
     sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output := sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_DUPLICATE_20ea LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_DUPLICATE_20ea_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2272_l2267_DUPLICATE_2f87 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2272_l2267_DUPLICATE_2f87_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_2674_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_8ba0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_f905_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_860e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_5867_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_DUPLICATE_20ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_DUPLICATE_20ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_DUPLICATE_20ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2272_l2264_l2279_l2267_DUPLICATE_7116_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2279_DUPLICATE_2ee7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_edcc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2259_l2264_l2279_l2267_DUPLICATE_e491_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2272_l2267_DUPLICATE_2f87_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2272_l2267_DUPLICATE_2f87_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2259_l2272_l2264_l2267_DUPLICATE_2bf6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_3fda_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2259_c1_b977] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2279_c7_4a47] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2279_c7_4a47] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2279_c7_4a47] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2279_c7_4a47] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;

     -- t8_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     t8_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     t8_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_b977_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_4a47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- printf_uxn_opcodes_h_l2260_c3_d844[uxn_opcodes_h_l2260_c3_d844] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2260_c3_d844_uxn_opcodes_h_l2260_c3_d844_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- t8_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     t8_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     t8_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2272_c7_58e3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_58e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2267_c7_1128] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;

     -- t8_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_1128_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2264_c7_535f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_535f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2259_c2_fdff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_12f7_uxn_opcodes_h_l2286_l2255_DUPLICATE_90ee LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_12f7_uxn_opcodes_h_l2286_l2255_DUPLICATE_90ee_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_12f7(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_fdff_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_12f7_uxn_opcodes_h_l2286_l2255_DUPLICATE_90ee_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_12f7_uxn_opcodes_h_l2286_l2255_DUPLICATE_90ee_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
