-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity neq_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_85d5529e;
architecture arch of neq_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1180_c6_76ef]
signal BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1180_c1_6b47]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1180_c2_be97]
signal n8_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1180_c2_be97]
signal t8_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1180_c2_be97]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1180_c2_be97]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1180_c2_be97]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1180_c2_be97]
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1180_c2_be97]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1180_c2_be97]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1181_c3_8ac6[uxn_opcodes_h_l1181_c3_8ac6]
signal printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1185_c11_09c3]
signal BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1185_c7_862c]
signal n8_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1185_c7_862c]
signal t8_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1185_c7_862c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1185_c7_862c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1185_c7_862c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1185_c7_862c]
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1185_c7_862c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1185_c7_862c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1188_c11_56d3]
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal n8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal t8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c7_dff7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1191_c11_ae6d]
signal BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal n8_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1191_c7_5e00]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1194_c30_d400]
signal sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1197_c21_f84c]
signal BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1197_c21_aae3]
signal MUX_uxn_opcodes_h_l1197_c21_aae3_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1197_c21_aae3_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1197_c21_aae3_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1197_c21_aae3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_b654]
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_96c6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_96c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_96c6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_left,
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_right,
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output);

-- n8_MUX_uxn_opcodes_h_l1180_c2_be97
n8_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
n8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
n8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- t8_MUX_uxn_opcodes_h_l1180_c2_be97
t8_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
t8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
t8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97
result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

-- printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6
printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6 : entity work.printf_uxn_opcodes_h_l1181_c3_8ac6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3
BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_left,
BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_right,
BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output);

-- n8_MUX_uxn_opcodes_h_l1185_c7_862c
n8_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
n8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
n8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- t8_MUX_uxn_opcodes_h_l1185_c7_862c
t8_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
t8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
t8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c
result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c
result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3
BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_left,
BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_right,
BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output);

-- n8_MUX_uxn_opcodes_h_l1188_c7_dff7
n8_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- t8_MUX_uxn_opcodes_h_l1188_c7_dff7
t8_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7
result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d
BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_left,
BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_right,
BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output);

-- n8_MUX_uxn_opcodes_h_l1191_c7_5e00
n8_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00
result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00
result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00
result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00
result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00
result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1194_c30_d400
sp_relative_shift_uxn_opcodes_h_l1194_c30_d400 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_ins,
sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_x,
sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_y,
sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c
BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_left,
BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_right,
BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output);

-- MUX_uxn_opcodes_h_l1197_c21_aae3
MUX_uxn_opcodes_h_l1197_c21_aae3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1197_c21_aae3_cond,
MUX_uxn_opcodes_h_l1197_c21_aae3_iftrue,
MUX_uxn_opcodes_h_l1197_c21_aae3_iffalse,
MUX_uxn_opcodes_h_l1197_c21_aae3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_left,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_right,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output,
 n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output,
 n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output,
 n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output,
 n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output,
 sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output,
 MUX_uxn_opcodes_h_l1197_c21_aae3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1182_c3_f1ea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_079b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1196_c3_c898 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1188_l1191_DUPLICATE_a204_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1176_l1205_DUPLICATE_59d7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_079b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_079b;
     VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1196_c3_c898 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1196_c3_c898;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1182_c3_f1ea := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1182_c3_f1ea;
     VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_iftrue := resize(to_unsigned(0, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1188_c11_56d3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1185_c11_09c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1191_c11_ae6d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1194_c30_d400] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_ins;
     sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_x;
     sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output := sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1197_c21_f84c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_b654] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_left;
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output := BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1188_l1191_DUPLICATE_a204 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1188_l1191_DUPLICATE_a204_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1180_c6_76ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_left;
     BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output := BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_76ef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1185_c11_09c3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c11_56d3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1191_c11_ae6d_return_output;
     VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1197_c21_f84c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_b654_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_fa4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1191_DUPLICATE_201d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_76a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1185_l1199_l1188_l1180_DUPLICATE_c6c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1188_l1191_DUPLICATE_a204_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1188_l1191_DUPLICATE_a204_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1185_l1188_l1180_l1191_DUPLICATE_e167_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1194_c30_d400_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_96c6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_96c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output;

     -- MUX[uxn_opcodes_h_l1197_c21_aae3] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1197_c21_aae3_cond <= VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_cond;
     MUX_uxn_opcodes_h_l1197_c21_aae3_iftrue <= VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_iftrue;
     MUX_uxn_opcodes_h_l1197_c21_aae3_iffalse <= VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_return_output := MUX_uxn_opcodes_h_l1197_c21_aae3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- n8_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1180_c1_6b47] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output;

     -- t8_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_96c6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue := VAR_MUX_uxn_opcodes_h_l1197_c21_aae3_return_output;
     VAR_printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1180_c1_6b47_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_96c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- printf_uxn_opcodes_h_l1181_c3_8ac6[uxn_opcodes_h_l1181_c3_8ac6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1181_c3_8ac6_uxn_opcodes_h_l1181_c3_8ac6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- t8_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     t8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     t8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- n8_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1191_c7_5e00] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1191_c7_5e00_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     n8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     n8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     t8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     t8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c7_dff7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c7_dff7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;
     -- n8_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     n8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     n8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1185_c7_862c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1185_c7_862c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1180_c2_be97] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1176_l1205_DUPLICATE_59d7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1176_l1205_DUPLICATE_59d7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_be97_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1180_c2_be97_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1176_l1205_DUPLICATE_59d7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1176_l1205_DUPLICATE_59d7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
