-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity sth_0CLK_d6c995e8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_d6c995e8;
architecture arch of sth_0CLK_d6c995e8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2601_c6_cf1c]
signal BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2601_c1_e30b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : signed(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2601_c2_9dbf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2602_c3_837a[uxn_opcodes_h_l2602_c3_837a]
signal printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2606_c11_ed35]
signal BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : signed(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2606_c7_4e4f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2609_c11_2fa1]
signal BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2609_c7_818f]
signal t8_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : signed(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2609_c7_818f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2612_c32_0acf]
signal BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2612_c32_6cd5]
signal BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2612_c32_96f3]
signal MUX_uxn_opcodes_h_l2612_c32_96f3_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2612_c32_96f3_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2612_c32_96f3_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2612_c32_96f3_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2614_c11_cda0]
signal BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : signed(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2614_c7_4867]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2618_c11_9c89]
signal BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2618_c7_1b87]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2618_c7_1b87]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2618_c7_1b87]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2618_c7_1b87]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2618_c7_1b87]
signal result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2618_c7_1b87]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_f6b2]
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2624_c7_8178]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_8178]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_8178]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_6621( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.stack_value := ref_toks_6;
      base.is_opc_done := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c
BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_left,
BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_right,
BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output);

-- t8_MUX_uxn_opcodes_h_l2601_c2_9dbf
t8_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf
result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

-- printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a
printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a : entity work.printf_uxn_opcodes_h_l2602_c3_837a_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35
BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_left,
BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_right,
BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output);

-- t8_MUX_uxn_opcodes_h_l2606_c7_4e4f
t8_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f
result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_left,
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_right,
BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output);

-- t8_MUX_uxn_opcodes_h_l2609_c7_818f
t8_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
t8_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
t8_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f
result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f
result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf
BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_left,
BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_right,
BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5
BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_left,
BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_right,
BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output);

-- MUX_uxn_opcodes_h_l2612_c32_96f3
MUX_uxn_opcodes_h_l2612_c32_96f3 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2612_c32_96f3_cond,
MUX_uxn_opcodes_h_l2612_c32_96f3_iftrue,
MUX_uxn_opcodes_h_l2612_c32_96f3_iffalse,
MUX_uxn_opcodes_h_l2612_c32_96f3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_left,
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_right,
BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867
result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_left,
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_right,
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87
result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87
result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_cond,
result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_left,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_right,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output,
 t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output,
 t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output,
 t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output,
 MUX_uxn_opcodes_h_l2612_c32_96f3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2603_c3_7e7b : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2607_c3_d29e : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2616_c3_7946 : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_b1d2 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2606_l2601_l2614_DUPLICATE_b5fd_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2618_l2609_l2614_DUPLICATE_9e90_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6621_uxn_opcodes_h_l2597_l2630_DUPLICATE_180d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2607_c3_d29e := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2607_c3_d29e;
     VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_right := to_unsigned(5, 3);
     VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_iffalse := resize(to_signed(-1, 2), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_b1d2 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_b1d2;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2616_c3_7946 := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2616_c3_7946;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_right := to_unsigned(128, 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2603_c3_7e7b := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2603_c3_7e7b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2606_c11_ed35] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_left;
     BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output := BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2606_l2601_l2614_DUPLICATE_b5fd LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2606_l2601_l2614_DUPLICATE_b5fd_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2618_l2609_l2614_DUPLICATE_9e90 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2618_l2609_l2614_DUPLICATE_9e90_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2614_c11_cda0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_f6b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2609_c11_2fa1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2601_c6_cf1c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2618_c11_9c89] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_left;
     BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output := BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2612_c32_0acf] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_left;
     BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output := BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2612_c32_0acf_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2601_c6_cf1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2606_c11_ed35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2609_c11_2fa1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2614_c11_cda0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_9c89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_f6b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2606_l2601_l2614_DUPLICATE_b5fd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2606_l2601_l2614_DUPLICATE_b5fd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2606_l2601_l2614_DUPLICATE_b5fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2609_l2606_l2624_l2618_l2614_DUPLICATE_32fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2606_l2618_l2601_l2614_DUPLICATE_5bb5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2618_DUPLICATE_9761_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2624_l2614_DUPLICATE_38d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2618_l2609_l2614_DUPLICATE_9e90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2618_l2609_l2614_DUPLICATE_9e90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2618_l2609_l2614_DUPLICATE_9e90_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2609_l2606_l2601_l2618_l2614_DUPLICATE_46a1_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_8178] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2601_c1_e30b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2618_c7_1b87] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2618_c7_1b87] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2624_c7_8178] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output;

     -- t8_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     t8_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     t8_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2612_c32_6cd5] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_left;
     BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output := BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_8178] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2618_c7_1b87] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output := result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2612_c32_6cd5_return_output;
     VAR_printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2601_c1_e30b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_8178_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2624_c7_8178_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_8178_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2618_c7_1b87] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- MUX[uxn_opcodes_h_l2612_c32_96f3] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2612_c32_96f3_cond <= VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_cond;
     MUX_uxn_opcodes_h_l2612_c32_96f3_iftrue <= VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_iftrue;
     MUX_uxn_opcodes_h_l2612_c32_96f3_iffalse <= VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_return_output := MUX_uxn_opcodes_h_l2612_c32_96f3_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2618_c7_1b87] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2618_c7_1b87] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;

     -- printf_uxn_opcodes_h_l2602_c3_837a[uxn_opcodes_h_l2602_c3_837a] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2602_c3_837a_uxn_opcodes_h_l2602_c3_837a_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue := VAR_MUX_uxn_opcodes_h_l2612_c32_96f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_1b87_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2614_c7_4867] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2614_c7_4867_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2609_c7_818f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2609_c7_818f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2606_c7_4e4f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2606_c7_4e4f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2601_c2_9dbf] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_6621_uxn_opcodes_h_l2597_l2630_DUPLICATE_180d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6621_uxn_opcodes_h_l2597_l2630_DUPLICATE_180d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_6621(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2601_c2_9dbf_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6621_uxn_opcodes_h_l2597_l2630_DUPLICATE_180d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6621_uxn_opcodes_h_l2597_l2630_DUPLICATE_180d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
