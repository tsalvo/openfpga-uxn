-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity equ_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_6d7675a8;
architecture arch of equ_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1226_c6_e17c]
signal BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1226_c1_d432]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1226_c2_524a]
signal n8_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1226_c2_524a]
signal t8_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1226_c2_524a]
signal result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1226_c2_524a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1226_c2_524a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1226_c2_524a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1226_c2_524a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1226_c2_524a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l1227_c3_9976[uxn_opcodes_h_l1227_c3_9976]
signal printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1231_c11_9f31]
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1231_c7_1ef5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1234_c11_3f43]
signal BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal n8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal t8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1234_c7_c71a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1238_c11_843a]
signal BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1238_c7_06df]
signal n8_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1238_c7_06df]
signal result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1238_c7_06df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1238_c7_06df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1238_c7_06df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1238_c7_06df]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1238_c7_06df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1241_c11_d127]
signal BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal n8_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1241_c7_7c62]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1244_c30_b982]
signal sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1247_c21_4306]
signal BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1247_c21_ee11]
signal MUX_uxn_opcodes_h_l1247_c21_ee11_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1247_c21_ee11_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1247_c21_ee11_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1247_c21_ee11_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1249_c11_3ae8]
signal BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1249_c7_3751]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1249_c7_3751]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1249_c7_3751]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c
BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_left,
BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_right,
BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output);

-- n8_MUX_uxn_opcodes_h_l1226_c2_524a
n8_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
n8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
n8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- t8_MUX_uxn_opcodes_h_l1226_c2_524a
t8_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
t8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
t8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a
result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a
result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a
result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a
result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

-- printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976
printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976 : entity work.printf_uxn_opcodes_h_l1227_c3_9976_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_left,
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_right,
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output);

-- n8_MUX_uxn_opcodes_h_l1231_c7_1ef5
n8_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- t8_MUX_uxn_opcodes_h_l1231_c7_1ef5
t8_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_left,
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_right,
BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output);

-- n8_MUX_uxn_opcodes_h_l1234_c7_c71a
n8_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- t8_MUX_uxn_opcodes_h_l1234_c7_c71a
t8_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a
BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_left,
BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_right,
BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output);

-- n8_MUX_uxn_opcodes_h_l1238_c7_06df
n8_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
n8_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
n8_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df
result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df
result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df
result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df
result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df
result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_left,
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_right,
BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output);

-- n8_MUX_uxn_opcodes_h_l1241_c7_7c62
n8_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1244_c30_b982
sp_relative_shift_uxn_opcodes_h_l1244_c30_b982 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_ins,
sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_x,
sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_y,
sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306
BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_left,
BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_right,
BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output);

-- MUX_uxn_opcodes_h_l1247_c21_ee11
MUX_uxn_opcodes_h_l1247_c21_ee11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1247_c21_ee11_cond,
MUX_uxn_opcodes_h_l1247_c21_ee11_iftrue,
MUX_uxn_opcodes_h_l1247_c21_ee11_iffalse,
MUX_uxn_opcodes_h_l1247_c21_ee11_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8
BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_left,
BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_right,
BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751
result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751
result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751
result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output,
 n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output,
 n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output,
 n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output,
 n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output,
 n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output,
 sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output,
 MUX_uxn_opcodes_h_l1247_c21_ee11_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1228_c3_eb61 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1232_c3_f153 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1236_c3_8b03 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1239_c3_1412 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1246_c3_2d0a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1241_c7_7c62_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1255_l1222_DUPLICATE_64c1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1228_c3_eb61 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1228_c3_eb61;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1239_c3_1412 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1239_c3_1412;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1236_c3_8b03 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1236_c3_8b03;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1246_c3_2d0a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1246_c3_2d0a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1232_c3_f153 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1232_c3_f153;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_iffalse := resize(to_unsigned(0, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1231_c11_9f31] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_left;
     BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output := BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1241_c11_d127] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_left;
     BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output := BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1234_c11_3f43] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_left;
     BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output := BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1241_c7_7c62_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1247_c21_4306] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_left;
     BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output := BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1244_c30_b982] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_ins;
     sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_x;
     sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output := sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1249_c11_3ae8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1238_c11_843a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1226_c6_e17c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output := result.u8_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1226_c6_e17c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_9f31_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1234_c11_3f43_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1238_c11_843a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1241_c11_d127_return_output;
     VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c21_4306_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1249_c11_3ae8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_044c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1249_l1241_l1238_l1234_l1231_DUPLICATE_219b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_0414_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1249_l1238_l1234_l1231_l1226_DUPLICATE_bf7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1241_l1238_l1234_l1231_l1226_DUPLICATE_d027_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1244_c30_b982_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- n8_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- MUX[uxn_opcodes_h_l1247_c21_ee11] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1247_c21_ee11_cond <= VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_cond;
     MUX_uxn_opcodes_h_l1247_c21_ee11_iftrue <= VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_iftrue;
     MUX_uxn_opcodes_h_l1247_c21_ee11_iffalse <= VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_return_output := MUX_uxn_opcodes_h_l1247_c21_ee11_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- t8_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1249_c7_3751] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1226_c1_d432] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1249_c7_3751] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1249_c7_3751] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue := VAR_MUX_uxn_opcodes_h_l1247_c21_ee11_return_output;
     VAR_printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1226_c1_d432_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1249_c7_3751_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1249_c7_3751_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1249_c7_3751_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- printf_uxn_opcodes_h_l1227_c3_9976[uxn_opcodes_h_l1227_c3_9976] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1227_c3_9976_uxn_opcodes_h_l1227_c3_9976_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     n8_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     n8_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1241_c7_7c62] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1241_c7_7c62_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     t8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     t8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1238_c7_06df] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1238_c7_06df_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;
     -- n8_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1234_c7_c71a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1234_c7_c71a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     n8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     n8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1231_c7_1ef5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_1ef5_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1226_c2_524a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1255_l1222_DUPLICATE_64c1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1255_l1222_DUPLICATE_64c1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1226_c2_524a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1226_c2_524a_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1255_l1222_DUPLICATE_64c1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1255_l1222_DUPLICATE_64c1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
