-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity neq_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_6d7675a8;
architecture arch of neq_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1314_c6_717a]
signal BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1314_c1_bf57]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal n8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1314_c2_7e09]
signal t8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1315_c3_0d76[uxn_opcodes_h_l1315_c3_0d76]
signal printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1319_c11_3c89]
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1319_c7_3155]
signal n8_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1319_c7_3155]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1319_c7_3155]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1319_c7_3155]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1319_c7_3155]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1319_c7_3155]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1319_c7_3155]
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1319_c7_3155]
signal t8_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1322_c11_599d]
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal n8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1322_c7_78ba]
signal t8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1326_c11_a9f3]
signal BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1326_c7_001c]
signal n8_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1326_c7_001c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1326_c7_001c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1326_c7_001c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1326_c7_001c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1326_c7_001c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1326_c7_001c]
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1329_c11_6098]
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal n8_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1329_c7_30d4]
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1332_c30_f504]
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1335_c21_2c98]
signal BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1335_c21_33ae]
signal MUX_uxn_opcodes_h_l1335_c21_33ae_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1335_c21_33ae_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1335_c21_33ae_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1335_c21_33ae_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1337_c11_325f]
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1337_c7_d2de]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1337_c7_d2de]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1337_c7_d2de]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_left,
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_right,
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output);

-- n8_MUX_uxn_opcodes_h_l1314_c2_7e09
n8_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- t8_MUX_uxn_opcodes_h_l1314_c2_7e09
t8_MUX_uxn_opcodes_h_l1314_c2_7e09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond,
t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue,
t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse,
t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

-- printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76
printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76 : entity work.printf_uxn_opcodes_h_l1315_c3_0d76_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_left,
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_right,
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output);

-- n8_MUX_uxn_opcodes_h_l1319_c7_3155
n8_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
n8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
n8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- t8_MUX_uxn_opcodes_h_l1319_c7_3155
t8_MUX_uxn_opcodes_h_l1319_c7_3155 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1319_c7_3155_cond,
t8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue,
t8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse,
t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_left,
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_right,
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output);

-- n8_MUX_uxn_opcodes_h_l1322_c7_78ba
n8_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- t8_MUX_uxn_opcodes_h_l1322_c7_78ba
t8_MUX_uxn_opcodes_h_l1322_c7_78ba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond,
t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue,
t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse,
t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_left,
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_right,
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output);

-- n8_MUX_uxn_opcodes_h_l1326_c7_001c
n8_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
n8_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
n8_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_left,
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_right,
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output);

-- n8_MUX_uxn_opcodes_h_l1329_c7_30d4
n8_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1332_c30_f504
sp_relative_shift_uxn_opcodes_h_l1332_c30_f504 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_ins,
sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_x,
sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_y,
sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_left,
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_right,
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output);

-- MUX_uxn_opcodes_h_l1335_c21_33ae
MUX_uxn_opcodes_h_l1335_c21_33ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1335_c21_33ae_cond,
MUX_uxn_opcodes_h_l1335_c21_33ae_iftrue,
MUX_uxn_opcodes_h_l1335_c21_33ae_iffalse,
MUX_uxn_opcodes_h_l1335_c21_33ae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_left,
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_right,
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output,
 n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output,
 n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output,
 n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output,
 n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output,
 n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output,
 sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output,
 MUX_uxn_opcodes_h_l1335_c21_33ae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1316_c3_64e1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1320_c3_2886 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1324_c3_fd50 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_9fbd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1334_c3_34c7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1329_c7_30d4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1343_l1310_DUPLICATE_d415_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1320_c3_2886 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1320_c3_2886;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_right := to_unsigned(5, 3);
     VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1334_c3_34c7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1334_c3_34c7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_9fbd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_9fbd;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1316_c3_64e1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1316_c3_64e1;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1324_c3_fd50 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1324_c3_fd50;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1326_c11_a9f3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1319_c11_3c89] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_left;
     BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output := BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1335_c21_2c98] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_left;
     BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output := BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1322_c11_599d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1329_c7_30d4_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1337_c11_325f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1314_c6_717a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1329_c11_6098] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_left;
     BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output := BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1332_c30_f504] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_ins;
     sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_x;
     sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output := sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_717a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_3c89_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_599d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_a9f3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_6098_return_output;
     VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2c98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_325f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_6e5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1337_DUPLICATE_f306_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_4ece_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1326_l1322_l1319_l1314_l1337_DUPLICATE_b9dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_15e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_f504_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1314_c1_bf57] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output;

     -- MUX[uxn_opcodes_h_l1335_c21_33ae] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1335_c21_33ae_cond <= VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_cond;
     MUX_uxn_opcodes_h_l1335_c21_33ae_iftrue <= VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_iftrue;
     MUX_uxn_opcodes_h_l1335_c21_33ae_iffalse <= VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_return_output := MUX_uxn_opcodes_h_l1335_c21_33ae_return_output;

     -- n8_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1337_c7_d2de] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output;

     -- t8_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1337_c7_d2de] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1337_c7_d2de] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue := VAR_MUX_uxn_opcodes_h_l1335_c21_33ae_return_output;
     VAR_printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_bf57_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_d2de_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- printf_uxn_opcodes_h_l1315_c3_0d76[uxn_opcodes_h_l1315_c3_0d76] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1315_c3_0d76_uxn_opcodes_h_l1315_c3_0d76_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     t8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     t8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     n8_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     n8_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1329_c7_30d4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_30d4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1326_c7_001c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_001c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;
     -- n8_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     n8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     n8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1322_c7_78ba] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output := result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_78ba_return_output;
     -- n8_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1319_c7_3155] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_3155_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1314_c2_7e09] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1343_l1310_DUPLICATE_d415 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1343_l1310_DUPLICATE_d415_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_7e09_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1343_l1310_DUPLICATE_d415_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1343_l1310_DUPLICATE_d415_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
