-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub1_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub1_0CLK_64d180f1;
architecture arch of sub1_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2461_c6_eb32]
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal n8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2461_c2_8be1]
signal t8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2474_c11_46d1]
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal n8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2474_c7_ad89]
signal t8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2477_c11_4fef]
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal n8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2477_c7_b2af]
signal t8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2480_c11_7623]
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2480_c7_a1dc]
signal n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2480_c7_a1dc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2480_c7_a1dc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2480_c7_a1dc]
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2480_c7_a1dc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2480_c7_a1dc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2482_c30_1a7f]
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2485_c21_f5d4]
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_left,
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_right,
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output);

-- n8_MUX_uxn_opcodes_h_l2461_c2_8be1
n8_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- t8_MUX_uxn_opcodes_h_l2461_c2_8be1
t8_MUX_uxn_opcodes_h_l2461_c2_8be1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond,
t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue,
t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse,
t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_left,
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_right,
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output);

-- n8_MUX_uxn_opcodes_h_l2474_c7_ad89
n8_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- t8_MUX_uxn_opcodes_h_l2474_c7_ad89
t8_MUX_uxn_opcodes_h_l2474_c7_ad89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond,
t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue,
t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse,
t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_left,
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_right,
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output);

-- n8_MUX_uxn_opcodes_h_l2477_c7_b2af
n8_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- t8_MUX_uxn_opcodes_h_l2477_c7_b2af
t8_MUX_uxn_opcodes_h_l2477_c7_b2af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond,
t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue,
t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse,
t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_left,
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_right,
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output);

-- n8_MUX_uxn_opcodes_h_l2480_c7_a1dc
n8_MUX_uxn_opcodes_h_l2480_c7_a1dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond,
n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue,
n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse,
n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_ins,
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_x,
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_y,
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_left,
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_right,
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output,
 n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output,
 n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output,
 n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output,
 n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output,
 sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_c42b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_455d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_90f3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_f403 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f6d9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_b92d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f1db_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_16e5_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2489_l2457_DUPLICATE_2131_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_455d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_455d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_f403 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_f403;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_90f3 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_90f3;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_c42b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_c42b;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2477_c11_4fef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_left;
     BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output := BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2474_c11_46d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_b92d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_b92d_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f1db LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f1db_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2480_c11_7623] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_left;
     BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output := BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2482_c30_1a7f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_ins;
     sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_x;
     sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output := sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2485_c21_f5d4] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2461_c6_eb32] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_left;
     BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output := BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f6d9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f6d9_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_16e5 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_16e5_return_output := result.stack_address_sp_offset;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529_return_output := result.u8_value;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_eb32_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_46d1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_4fef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7623_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_f5d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f6d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f6d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f6d9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f1db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f1db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_f1db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_b92d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_b92d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_b92d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_16e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_16e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_2529_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_8be1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a7f_return_output;
     -- t8_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2480_c7_a1dc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2480_c7_a1dc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;

     -- n8_MUX[uxn_opcodes_h_l2480_c7_a1dc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond;
     n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue;
     n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output := n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2480_c7_a1dc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2480_c7_a1dc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2480_c7_a1dc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_a1dc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     -- t8_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- n8_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2477_c7_b2af] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_b2af_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- n8_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- t8_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2474_c7_ad89] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output := result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ad89_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- n8_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2461_c2_8be1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2489_l2457_DUPLICATE_2131 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2489_l2457_DUPLICATE_2131_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_8be1_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2489_l2457_DUPLICATE_2131_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2489_l2457_DUPLICATE_2131_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
