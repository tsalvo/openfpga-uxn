-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity jmp2_0CLK_9101a1df is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_9101a1df;
architecture arch of jmp2_0CLK_9101a1df is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l652_c6_b97f]
signal BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l652_c1_404d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l652_c2_bf08]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l652_c2_bf08]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l652_c2_bf08]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l652_c2_bf08]
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l652_c2_bf08]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l652_c2_bf08]
signal result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l652_c2_bf08]
signal t16_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l653_c3_78dc[uxn_opcodes_h_l653_c3_78dc]
signal printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l657_c11_cd53]
signal BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l657_c7_e218]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l657_c7_e218]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l657_c7_e218]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l657_c7_e218]
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l657_c7_e218]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l657_c7_e218]
signal result_pc_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l657_c7_e218]
signal t16_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l660_c11_e438]
signal BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l660_c7_5014]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l660_c7_5014]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l660_c7_5014]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l660_c7_5014]
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l660_c7_5014]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l660_c7_5014]
signal result_pc_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l660_c7_5014]
signal t16_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l662_c3_1b08]
signal CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l665_c11_822f]
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l665_c7_2d1a]
signal t16_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l668_c11_fe9d]
signal BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l668_c7_9566]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l668_c7_9566]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l668_c7_9566]
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l668_c7_9566]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l668_c7_9566]
signal result_pc_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l668_c7_9566]
signal t16_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l669_c3_931a]
signal BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output : unsigned(15 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l671_c32_56f1]
signal BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l671_c32_bc4f]
signal BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l671_c32_0776]
signal MUX_uxn_opcodes_h_l671_c32_0776_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l671_c32_0776_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l671_c32_0776_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l671_c32_0776_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l675_c11_67e9]
signal BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l675_c7_c417]
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l675_c7_c417]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l675_c7_c417]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_af99( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_pc_updated := ref_toks_5;
      base.pc := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f
BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_left,
BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_right,
BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- result_pc_MUX_uxn_opcodes_h_l652_c2_bf08
result_pc_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- t16_MUX_uxn_opcodes_h_l652_c2_bf08
t16_MUX_uxn_opcodes_h_l652_c2_bf08 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l652_c2_bf08_cond,
t16_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue,
t16_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse,
t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

-- printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc
printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc : entity work.printf_uxn_opcodes_h_l653_c3_78dc_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53
BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_left,
BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_right,
BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- result_pc_MUX_uxn_opcodes_h_l657_c7_e218
result_pc_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l657_c7_e218_cond,
result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- t16_MUX_uxn_opcodes_h_l657_c7_e218
t16_MUX_uxn_opcodes_h_l657_c7_e218 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l657_c7_e218_cond,
t16_MUX_uxn_opcodes_h_l657_c7_e218_iftrue,
t16_MUX_uxn_opcodes_h_l657_c7_e218_iffalse,
t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438
BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_left,
BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_right,
BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- result_pc_MUX_uxn_opcodes_h_l660_c7_5014
result_pc_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l660_c7_5014_cond,
result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- t16_MUX_uxn_opcodes_h_l660_c7_5014
t16_MUX_uxn_opcodes_h_l660_c7_5014 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l660_c7_5014_cond,
t16_MUX_uxn_opcodes_h_l660_c7_5014_iftrue,
t16_MUX_uxn_opcodes_h_l660_c7_5014_iffalse,
t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output);

-- CONST_SL_8_uxn_opcodes_h_l662_c3_1b08
CONST_SL_8_uxn_opcodes_h_l662_c3_1b08 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_x,
CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f
BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_left,
BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_right,
BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a
result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- t16_MUX_uxn_opcodes_h_l665_c7_2d1a
t16_MUX_uxn_opcodes_h_l665_c7_2d1a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l665_c7_2d1a_cond,
t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue,
t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse,
t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d
BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_left,
BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_right,
BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output);

-- result_pc_MUX_uxn_opcodes_h_l668_c7_9566
result_pc_MUX_uxn_opcodes_h_l668_c7_9566 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l668_c7_9566_cond,
result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iftrue,
result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iffalse,
result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output);

-- t16_MUX_uxn_opcodes_h_l668_c7_9566
t16_MUX_uxn_opcodes_h_l668_c7_9566 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l668_c7_9566_cond,
t16_MUX_uxn_opcodes_h_l668_c7_9566_iftrue,
t16_MUX_uxn_opcodes_h_l668_c7_9566_iffalse,
t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l669_c3_931a
BIN_OP_OR_uxn_opcodes_h_l669_c3_931a : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_left,
BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_right,
BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1
BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_left,
BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_right,
BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f
BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_left,
BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_right,
BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output);

-- MUX_uxn_opcodes_h_l671_c32_0776
MUX_uxn_opcodes_h_l671_c32_0776 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l671_c32_0776_cond,
MUX_uxn_opcodes_h_l671_c32_0776_iftrue,
MUX_uxn_opcodes_h_l671_c32_0776_iffalse,
MUX_uxn_opcodes_h_l671_c32_0776_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9
BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_left,
BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_right,
BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output,
 CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output,
 result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output,
 t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output,
 BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output,
 BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output,
 BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output,
 MUX_uxn_opcodes_h_l671_c32_0776_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l654_c3_4671 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_765b : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l663_c3_069c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l666_c3_d447 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l665_c7_2d1a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l671_c32_0776_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l671_c32_0776_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l671_c32_0776_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l671_c32_0776_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l669_l661_DUPLICATE_329b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_af99_uxn_opcodes_h_l648_l681_DUPLICATE_5f10_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_right := to_unsigned(3, 2);
     VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l654_c3_4671 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l654_c3_4671;
     VAR_MUX_uxn_opcodes_h_l671_c32_0776_iffalse := resize(to_signed(-2, 3), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_765b := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_765b;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l666_c3_d447 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l666_c3_d447;
     VAR_MUX_uxn_opcodes_h_l671_c32_0776_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_right := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_right := to_unsigned(128, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l663_c3_069c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l663_c3_069c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_iffalse := t16;
     -- BIN_OP_AND[uxn_opcodes_h_l671_c32_56f1] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_left;
     BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output := BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l675_c11_67e9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_left;
     BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output := BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l665_c11_822f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_left;
     BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output := BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l660_c11_e438] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_left;
     BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output := BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l657_c11_cd53] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_left;
     BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output := BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output := result.pc;

     -- BIN_OP_EQ[uxn_opcodes_h_l668_c11_fe9d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_left;
     BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output := BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l652_c6_b97f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_left;
     BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output := BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l669_l661_DUPLICATE_329b LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l669_l661_DUPLICATE_329b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l665_c7_2d1a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_left := VAR_BIN_OP_AND_uxn_opcodes_h_l671_c32_56f1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_b97f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_cd53_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_e438_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_822f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_fe9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_67e9_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l669_l661_DUPLICATE_329b_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l669_l661_DUPLICATE_329b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_c31e_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_e2f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l675_l668_l657_DUPLICATE_1632_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_7502_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l675_l652_l657_DUPLICATE_482c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l665_c7_2d1a_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l652_c1_404d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l675_c7_c417] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l662_c3_1b08] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_x <= VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output := CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l675_c7_c417] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l675_c7_c417] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l669_c3_931a] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_left;
     BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output := BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l671_c32_bc4f] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_left;
     BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output := BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l671_c32_0776_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l671_c32_bc4f_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_931a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_1b08_return_output;
     VAR_printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l652_c1_404d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_c417_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_c417_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_c417_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l668_c7_9566] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l668_c7_9566] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l668_c7_9566_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_cond;
     result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iftrue;
     result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output := result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l668_c7_9566] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output;

     -- t16_MUX[uxn_opcodes_h_l668_c7_9566] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l668_c7_9566_cond <= VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_cond;
     t16_MUX_uxn_opcodes_h_l668_c7_9566_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_iftrue;
     t16_MUX_uxn_opcodes_h_l668_c7_9566_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output := t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l668_c7_9566] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output;

     -- printf_uxn_opcodes_h_l653_c3_78dc[uxn_opcodes_h_l653_c3_78dc] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l653_c3_78dc_uxn_opcodes_h_l653_c3_78dc_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- MUX[uxn_opcodes_h_l671_c32_0776] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l671_c32_0776_cond <= VAR_MUX_uxn_opcodes_h_l671_c32_0776_cond;
     MUX_uxn_opcodes_h_l671_c32_0776_iftrue <= VAR_MUX_uxn_opcodes_h_l671_c32_0776_iftrue;
     MUX_uxn_opcodes_h_l671_c32_0776_iffalse <= VAR_MUX_uxn_opcodes_h_l671_c32_0776_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l671_c32_0776_return_output := MUX_uxn_opcodes_h_l671_c32_0776_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue := VAR_MUX_uxn_opcodes_h_l671_c32_0776_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_9566_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_9566_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l668_c7_9566_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l668_c7_9566_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l668_c7_9566] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- t16_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_9566_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_t16_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l665_c7_2d1a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output := result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- t16_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     t16_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     t16_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output := t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_2d1a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_t16_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     -- t16_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     t16_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     t16_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output := t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l660_c7_5014] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output := result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_5014_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_t16_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     -- result_pc_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l657_c7_e218] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output;

     -- t16_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     t16_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     t16_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- Submodule level 7
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_e218_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l652_c2_bf08] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_af99_uxn_opcodes_h_l648_l681_DUPLICATE_5f10 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_af99_uxn_opcodes_h_l648_l681_DUPLICATE_5f10_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_af99(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_bf08_return_output,
     VAR_result_pc_MUX_uxn_opcodes_h_l652_c2_bf08_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_af99_uxn_opcodes_h_l648_l681_DUPLICATE_5f10_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_af99_uxn_opcodes_h_l648_l681_DUPLICATE_5f10_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
