-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity ldz_0CLK_df07acae is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_df07acae;
architecture arch of ldz_0CLK_df07acae is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1553_c6_7b41]
signal BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1553_c1_cac0]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal t8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(15 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1553_c2_41bc]
signal tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1554_c3_510b[uxn_opcodes_h_l1554_c3_510b]
signal printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1558_c11_9138]
signal BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal t8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(15 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1558_c7_cef5]
signal tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1561_c11_e7c7]
signal BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(15 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1561_c7_d5a4]
signal tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1564_c32_bf3a]
signal BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1564_c32_f035]
signal BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1564_c32_f737]
signal MUX_uxn_opcodes_h_l1564_c32_f737_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1564_c32_f737_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1564_c32_f737_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1564_c32_f737_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1567_c11_3643]
signal BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(15 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1567_c7_6c32]
signal tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1571_c11_4cf0]
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1571_c7_86b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1571_c7_86b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1571_c7_86b9]
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1571_c7_86b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1571_c7_86b9]
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1577_c11_9d7a]
signal BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1577_c7_9f6e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1577_c7_9f6e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_3413( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.ram_addr := ref_toks_6;
      base.stack_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41
BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_left,
BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_right,
BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output);

-- t8_MUX_uxn_opcodes_h_l1553_c2_41bc
t8_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc
result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc
result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc
result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc
result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc
result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc
tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond,
tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue,
tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse,
tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

-- printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b
printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b : entity work.printf_uxn_opcodes_h_l1554_c3_510b_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138
BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_left,
BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_right,
BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output);

-- t8_MUX_uxn_opcodes_h_l1558_c7_cef5
t8_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5
result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5
result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5
result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5
result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5
result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5
tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond,
tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue,
tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse,
tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7
BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_left,
BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_right,
BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output);

-- t8_MUX_uxn_opcodes_h_l1561_c7_d5a4
t8_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4
result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4
tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond,
tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue,
tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse,
tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a
BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_left,
BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_right,
BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035
BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_left,
BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_right,
BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output);

-- MUX_uxn_opcodes_h_l1564_c32_f737
MUX_uxn_opcodes_h_l1564_c32_f737 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1564_c32_f737_cond,
MUX_uxn_opcodes_h_l1564_c32_f737_iftrue,
MUX_uxn_opcodes_h_l1564_c32_f737_iffalse,
MUX_uxn_opcodes_h_l1564_c32_f737_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643
BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_left,
BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_right,
BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32
result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32
result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32
result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32
result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32
result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32
tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_cond,
tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue,
tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse,
tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_left,
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_right,
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_cond,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9
tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_cond,
tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue,
tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse,
tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_left,
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_right,
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e
result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output,
 t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output,
 t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output,
 t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output,
 MUX_uxn_opcodes_h_l1564_c32_f737_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output,
 tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1555_c3_faa7 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_6aa8 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1564_c32_f737_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1564_c32_f737_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1564_c32_f737_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1564_c32_f737_return_output : signed(7 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1565_c21_56c0_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_2dc4_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1574_c3_43f7 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1553_l1558_l1561_DUPLICATE_d57c_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_8790_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_f7f9_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1567_l1571_l1561_DUPLICATE_0b04_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3413_uxn_opcodes_h_l1582_l1549_DUPLICATE_b892_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_right := to_unsigned(3, 2);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1574_c3_43f7 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1574_c3_43f7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_6aa8 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_6aa8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1555_c3_faa7 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1555_c3_faa7;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1564_c32_f737_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1564_c32_f737_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_left := VAR_phase;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse := tmp8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1567_l1571_l1561_DUPLICATE_0b04 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1567_l1571_l1561_DUPLICATE_0b04_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_f7f9 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_f7f9_return_output := result.ram_addr;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_8790 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_8790_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1553_c6_7b41] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_left;
     BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output := BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1569_c21_2dc4] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_2dc4_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1577_c11_9d7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1571_c11_4cf0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1561_c11_e7c7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1565_c21_56c0] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1565_c21_56c0_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1558_c11_9138] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_left;
     BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output := BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1553_l1558_l1561_DUPLICATE_d57c LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1553_l1558_l1561_DUPLICATE_d57c_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1567_c11_3643] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_left;
     BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output := BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output := result.is_stack_write;

     -- BIN_OP_AND[uxn_opcodes_h_l1564_c32_bf3a] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_left;
     BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output := BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1564_c32_bf3a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1553_c6_7b41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1558_c11_9138_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1561_c11_e7c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1567_c11_3643_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_4cf0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_9d7a_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1565_c21_56c0_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_2dc4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1553_l1558_l1561_DUPLICATE_d57c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1553_l1558_l1561_DUPLICATE_d57c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1553_l1558_l1561_DUPLICATE_d57c_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_f7f9_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_f7f9_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_f7f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1567_l1558_l1577_l1571_l1561_DUPLICATE_18a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_8790_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_8790_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1567_l1553_l1558_DUPLICATE_8790_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1577_l1561_DUPLICATE_8eed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1567_l1571_l1561_DUPLICATE_0b04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1567_l1571_l1561_DUPLICATE_0b04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1567_l1571_l1561_DUPLICATE_0b04_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1567_l1553_l1558_l1571_l1561_DUPLICATE_c7ff_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- t8_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1571_c7_86b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1553_c1_cac0] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1564_c32_f035] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_left;
     BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output := BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1577_c7_9f6e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1571_c7_86b9] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output := result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1577_c7_9f6e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1571_c7_86b9] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_cond;
     tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output := tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1564_c32_f737_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1564_c32_f035_return_output;
     VAR_printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1553_c1_cac0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1577_c7_9f6e_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;
     -- MUX[uxn_opcodes_h_l1564_c32_f737] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1564_c32_f737_cond <= VAR_MUX_uxn_opcodes_h_l1564_c32_f737_cond;
     MUX_uxn_opcodes_h_l1564_c32_f737_iftrue <= VAR_MUX_uxn_opcodes_h_l1564_c32_f737_iftrue;
     MUX_uxn_opcodes_h_l1564_c32_f737_iffalse <= VAR_MUX_uxn_opcodes_h_l1564_c32_f737_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1564_c32_f737_return_output := MUX_uxn_opcodes_h_l1564_c32_f737_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1571_c7_86b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1571_c7_86b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- printf_uxn_opcodes_h_l1554_c3_510b[uxn_opcodes_h_l1554_c3_510b] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1554_c3_510b_uxn_opcodes_h_l1554_c3_510b_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue := VAR_MUX_uxn_opcodes_h_l1564_c32_f737_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_86b9_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1567_c7_6c32] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1567_c7_6c32_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1561_c7_d5a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1561_c7_d5a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1558_c7_cef5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1558_c7_cef5_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1553_c2_41bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3413_uxn_opcodes_h_l1582_l1549_DUPLICATE_b892 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3413_uxn_opcodes_h_l1582_l1549_DUPLICATE_b892_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3413(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1553_c2_41bc_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3413_uxn_opcodes_h_l1582_l1549_DUPLICATE_b892_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3413_uxn_opcodes_h_l1582_l1549_DUPLICATE_b892_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
