-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity jsr2_0CLK_609876da is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr2_0CLK_609876da;
architecture arch of jsr2_0CLK_609876da is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l774_c6_fc02]
signal BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l774_c2_9818]
signal t16_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l774_c2_9818]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l787_c11_6396]
signal BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l787_c7_00d4]
signal t16_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l787_c7_00d4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l790_c11_902d]
signal BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal t16_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l790_c7_2b5e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l792_c3_6568]
signal CONST_SL_8_uxn_opcodes_h_l792_c3_6568_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l793_c30_a693]
signal sp_relative_shift_uxn_opcodes_h_l793_c30_a693_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l793_c30_a693_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l793_c30_a693_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l795_c11_d02d]
signal BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal t16_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l795_c7_8f4a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l796_c3_87a0]
signal BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l803_c11_84c1]
signal BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l803_c7_edb3]
signal result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l803_c7_edb3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l803_c7_edb3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l803_c7_edb3]
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l803_c7_edb3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l803_c7_edb3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : signed(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l806_c31_1137]
signal CONST_SR_8_uxn_opcodes_h_l806_c31_1137_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output : unsigned(15 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_d9be( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.is_pc_updated := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.sp_relative_shift := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02
BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_left,
BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_right,
BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output);

-- t16_MUX_uxn_opcodes_h_l774_c2_9818
t16_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l774_c2_9818_cond,
t16_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
t16_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818
result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818
result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818
result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818
result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818
result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818
result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396
BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_left,
BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_right,
BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output);

-- t16_MUX_uxn_opcodes_h_l787_c7_00d4
t16_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
t16_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
t16_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4
result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4
result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4
result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4
result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4
result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4
result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d
BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_left,
BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_right,
BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output);

-- t16_MUX_uxn_opcodes_h_l790_c7_2b5e
t16_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e
result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e
result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e
result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e
result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e
result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output);

-- CONST_SL_8_uxn_opcodes_h_l792_c3_6568
CONST_SL_8_uxn_opcodes_h_l792_c3_6568 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l792_c3_6568_x,
CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output);

-- sp_relative_shift_uxn_opcodes_h_l793_c30_a693
sp_relative_shift_uxn_opcodes_h_l793_c30_a693 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l793_c30_a693_ins,
sp_relative_shift_uxn_opcodes_h_l793_c30_a693_x,
sp_relative_shift_uxn_opcodes_h_l793_c30_a693_y,
sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d
BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_left,
BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_right,
BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output);

-- t16_MUX_uxn_opcodes_h_l795_c7_8f4a
t16_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a
result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a
result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a
result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0
BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_left,
BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_right,
BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1
BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_left,
BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_right,
BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3
result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond,
result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3
result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3
result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond,
result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output);

-- CONST_SR_8_uxn_opcodes_h_l806_c31_1137
CONST_SR_8_uxn_opcodes_h_l806_c31_1137 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l806_c31_1137_x,
CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output,
 t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output,
 t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output,
 t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output,
 CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output,
 sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output,
 t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output,
 BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output,
 CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l784_c3_7960 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l779_c3_2b68 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l788_c3_40cc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l792_c3_6568_x : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l800_c3_a40b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l798_c3_10fb : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l801_c21_f6a0_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l805_c3_9826 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l804_c3_f37b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l806_c31_1137_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l806_c21_2be7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_2ae2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_0cc7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l787_l803_DUPLICATE_2ef9_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l796_l791_DUPLICATE_8800_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l803_l790_DUPLICATE_969c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l812_l770_DUPLICATE_47fb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l805_c3_9826 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l805_c3_9826;
     VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_right := to_unsigned(2, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l800_c3_a40b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l800_c3_a40b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l784_c3_7960 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l784_c3_7960;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l788_c3_40cc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l788_c3_40cc;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l804_c3_f37b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l804_c3_f37b;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l779_c3_2b68 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l779_c3_2b68;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_right := to_unsigned(4, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l798_c3_10fb := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l798_c3_10fb;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_ins := VAR_ins;
     VAR_CONST_SR_8_uxn_opcodes_h_l806_c31_1137_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_0cc7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_0cc7_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l803_c11_84c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_left;
     BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output := BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l774_c6_fc02] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_left;
     BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output := BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l774_c2_9818_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l787_l803_DUPLICATE_2ef9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l787_l803_DUPLICATE_2ef9_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l790_c11_902d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_left;
     BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output := BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3_return_output := result.u8_value;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output := result.u16_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l774_c2_9818_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l795_c11_d02d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_left;
     BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output := BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l801_c21_f6a0] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l801_c21_f6a0_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- sp_relative_shift[uxn_opcodes_h_l793_c30_a693] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l793_c30_a693_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_ins;
     sp_relative_shift_uxn_opcodes_h_l793_c30_a693_x <= VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_x;
     sp_relative_shift_uxn_opcodes_h_l793_c30_a693_y <= VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output := sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l787_c11_6396] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_left;
     BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output := BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l803_l790_DUPLICATE_969c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l803_l790_DUPLICATE_969c_return_output := result.stack_address_sp_offset;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l796_l791_DUPLICATE_8800 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l796_l791_DUPLICATE_8800_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_SR_8[uxn_opcodes_h_l806_c31_1137] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l806_c31_1137_x <= VAR_CONST_SR_8_uxn_opcodes_h_l806_c31_1137_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output := CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_2ae2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_2ae2_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c6_fc02_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l787_c11_6396_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l790_c11_902d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l795_c11_d02d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_84c1_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l796_l791_DUPLICATE_8800_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l792_c3_6568_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l796_l791_DUPLICATE_8800_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l801_c21_f6a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l787_l803_DUPLICATE_2ef9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l787_l803_DUPLICATE_2ef9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l790_l787_l774_l803_l795_DUPLICATE_a568_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_9fa8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l787_l803_l790_l795_DUPLICATE_db40_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_0cc7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_0cc7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_0cc7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_2ae2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_2ae2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l787_l790_l795_DUPLICATE_2ae2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l803_l790_DUPLICATE_969c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l803_l790_DUPLICATE_969c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l787_l803_l790_l774_DUPLICATE_37e3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l774_c2_9818_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l774_c2_9818_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l793_c30_a693_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l803_c7_edb3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l803_c7_edb3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l803_c7_edb3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l803_c7_edb3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l792_c3_6568] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l792_c3_6568_x <= VAR_CONST_SL_8_uxn_opcodes_h_l792_c3_6568_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output := CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l806_c21_2be7] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l806_c21_2be7_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l806_c31_1137_return_output);

     -- result_u16_value_MUX[uxn_opcodes_h_l803_c7_edb3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output := result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l796_c3_87a0] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_left;
     BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output := BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l796_c3_87a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l806_c21_2be7_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l792_c3_6568_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l803_c7_edb3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output := result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- t16_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_edb3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_t16_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- t16_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l795_c7_8f4a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output := result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l795_c7_8f4a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_t16_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l790_c7_2b5e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output := result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;

     -- t16_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     t16_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     t16_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l790_c7_2b5e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_t16_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l787_c7_00d4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output := result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- t16_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     t16_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     t16_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output := t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l787_c7_00d4_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l774_c2_9818_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l774_c2_9818] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_cond;
     result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output := result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l812_l770_DUPLICATE_47fb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l812_l770_DUPLICATE_47fb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d9be(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l774_c2_9818_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c2_9818_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l812_l770_DUPLICATE_47fb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l812_l770_DUPLICATE_47fb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
