-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 19
entity uint16_mux16_0CLK_4e6656cf is
port(
 sel : in unsigned(3 downto 0);
 in0 : in unsigned(15 downto 0);
 in1 : in unsigned(15 downto 0);
 in2 : in unsigned(15 downto 0);
 in3 : in unsigned(15 downto 0);
 in4 : in unsigned(15 downto 0);
 in5 : in unsigned(15 downto 0);
 in6 : in unsigned(15 downto 0);
 in7 : in unsigned(15 downto 0);
 in8 : in unsigned(15 downto 0);
 in9 : in unsigned(15 downto 0);
 in10 : in unsigned(15 downto 0);
 in11 : in unsigned(15 downto 0);
 in12 : in unsigned(15 downto 0);
 in13 : in unsigned(15 downto 0);
 in14 : in unsigned(15 downto 0);
 in15 : in unsigned(15 downto 0);
 return_output : out unsigned(15 downto 0));
end uint16_mux16_0CLK_4e6656cf;
architecture arch of uint16_mux16_0CLK_4e6656cf is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_8dfa]
signal layer0_node0_MUX_bit_math_h_l18_c3_8dfa_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iftrue : unsigned(15 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iffalse : unsigned(15 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output : unsigned(15 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_ee77]
signal layer0_node1_MUX_bit_math_h_l29_c3_ee77_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_ee77_iftrue : unsigned(15 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_ee77_iffalse : unsigned(15 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output : unsigned(15 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_55a7]
signal layer0_node2_MUX_bit_math_h_l40_c3_55a7_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_55a7_iftrue : unsigned(15 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_55a7_iffalse : unsigned(15 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output : unsigned(15 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_0c13]
signal layer0_node3_MUX_bit_math_h_l51_c3_0c13_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_0c13_iftrue : unsigned(15 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_0c13_iffalse : unsigned(15 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output : unsigned(15 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_ee64]
signal layer0_node4_MUX_bit_math_h_l62_c3_ee64_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_ee64_iftrue : unsigned(15 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_ee64_iffalse : unsigned(15 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output : unsigned(15 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_6697]
signal layer0_node5_MUX_bit_math_h_l73_c3_6697_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_6697_iftrue : unsigned(15 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_6697_iffalse : unsigned(15 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output : unsigned(15 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_d7ea]
signal layer0_node6_MUX_bit_math_h_l84_c3_d7ea_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iftrue : unsigned(15 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iffalse : unsigned(15 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output : unsigned(15 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_c417]
signal layer0_node7_MUX_bit_math_h_l95_c3_c417_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c417_iftrue : unsigned(15 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c417_iffalse : unsigned(15 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output : unsigned(15 downto 0);

-- layer1_node0_MUX[bit_math_h_l112_c3_a151]
signal layer1_node0_MUX_bit_math_h_l112_c3_a151_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_a151_iftrue : unsigned(15 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_a151_iffalse : unsigned(15 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output : unsigned(15 downto 0);

-- layer1_node1_MUX[bit_math_h_l123_c3_f7f1]
signal layer1_node1_MUX_bit_math_h_l123_c3_f7f1_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iftrue : unsigned(15 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iffalse : unsigned(15 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output : unsigned(15 downto 0);

-- layer1_node2_MUX[bit_math_h_l134_c3_5a40]
signal layer1_node2_MUX_bit_math_h_l134_c3_5a40_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_5a40_iftrue : unsigned(15 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_5a40_iffalse : unsigned(15 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output : unsigned(15 downto 0);

-- layer1_node3_MUX[bit_math_h_l145_c3_b458]
signal layer1_node3_MUX_bit_math_h_l145_c3_b458_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_b458_iftrue : unsigned(15 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_b458_iffalse : unsigned(15 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output : unsigned(15 downto 0);

-- layer2_node0_MUX[bit_math_h_l162_c3_9803]
signal layer2_node0_MUX_bit_math_h_l162_c3_9803_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_9803_iftrue : unsigned(15 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_9803_iffalse : unsigned(15 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output : unsigned(15 downto 0);

-- layer2_node1_MUX[bit_math_h_l173_c3_c834]
signal layer2_node1_MUX_bit_math_h_l173_c3_c834_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_c834_iftrue : unsigned(15 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_c834_iffalse : unsigned(15 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output : unsigned(15 downto 0);

-- layer3_node0_MUX[bit_math_h_l190_c3_d7d1]
signal layer3_node0_MUX_bit_math_h_l190_c3_d7d1_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iftrue : unsigned(15 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iffalse : unsigned(15 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output : unsigned(15 downto 0);

function uint4_0_0( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint4_1_1( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint4_2_2( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint4_3_3( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_8dfa
layer0_node0_MUX_bit_math_h_l18_c3_8dfa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_8dfa_cond,
layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_ee77
layer0_node1_MUX_bit_math_h_l29_c3_ee77 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_ee77_cond,
layer0_node1_MUX_bit_math_h_l29_c3_ee77_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_ee77_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_55a7
layer0_node2_MUX_bit_math_h_l40_c3_55a7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_55a7_cond,
layer0_node2_MUX_bit_math_h_l40_c3_55a7_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_55a7_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_0c13
layer0_node3_MUX_bit_math_h_l51_c3_0c13 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_0c13_cond,
layer0_node3_MUX_bit_math_h_l51_c3_0c13_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_0c13_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_ee64
layer0_node4_MUX_bit_math_h_l62_c3_ee64 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_ee64_cond,
layer0_node4_MUX_bit_math_h_l62_c3_ee64_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_ee64_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_6697
layer0_node5_MUX_bit_math_h_l73_c3_6697 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_6697_cond,
layer0_node5_MUX_bit_math_h_l73_c3_6697_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_6697_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_d7ea
layer0_node6_MUX_bit_math_h_l84_c3_d7ea : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_d7ea_cond,
layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_c417
layer0_node7_MUX_bit_math_h_l95_c3_c417 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_c417_cond,
layer0_node7_MUX_bit_math_h_l95_c3_c417_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_c417_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output);

-- layer1_node0_MUX_bit_math_h_l112_c3_a151
layer1_node0_MUX_bit_math_h_l112_c3_a151 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l112_c3_a151_cond,
layer1_node0_MUX_bit_math_h_l112_c3_a151_iftrue,
layer1_node0_MUX_bit_math_h_l112_c3_a151_iffalse,
layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output);

-- layer1_node1_MUX_bit_math_h_l123_c3_f7f1
layer1_node1_MUX_bit_math_h_l123_c3_f7f1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l123_c3_f7f1_cond,
layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iftrue,
layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iffalse,
layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output);

-- layer1_node2_MUX_bit_math_h_l134_c3_5a40
layer1_node2_MUX_bit_math_h_l134_c3_5a40 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l134_c3_5a40_cond,
layer1_node2_MUX_bit_math_h_l134_c3_5a40_iftrue,
layer1_node2_MUX_bit_math_h_l134_c3_5a40_iffalse,
layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output);

-- layer1_node3_MUX_bit_math_h_l145_c3_b458
layer1_node3_MUX_bit_math_h_l145_c3_b458 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l145_c3_b458_cond,
layer1_node3_MUX_bit_math_h_l145_c3_b458_iftrue,
layer1_node3_MUX_bit_math_h_l145_c3_b458_iffalse,
layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output);

-- layer2_node0_MUX_bit_math_h_l162_c3_9803
layer2_node0_MUX_bit_math_h_l162_c3_9803 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l162_c3_9803_cond,
layer2_node0_MUX_bit_math_h_l162_c3_9803_iftrue,
layer2_node0_MUX_bit_math_h_l162_c3_9803_iffalse,
layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output);

-- layer2_node1_MUX_bit_math_h_l173_c3_c834
layer2_node1_MUX_bit_math_h_l173_c3_c834 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l173_c3_c834_cond,
layer2_node1_MUX_bit_math_h_l173_c3_c834_iftrue,
layer2_node1_MUX_bit_math_h_l173_c3_c834_iffalse,
layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output);

-- layer3_node0_MUX_bit_math_h_l190_c3_d7d1
layer3_node0_MUX_bit_math_h_l190_c3_d7d1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l190_c3_d7d1_cond,
layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iftrue,
layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iffalse,
layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output,
 layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output,
 layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output,
 layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output,
 layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output,
 layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output,
 layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output,
 layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(15 downto 0);
 variable VAR_sel : unsigned(3 downto 0);
 variable VAR_in0 : unsigned(15 downto 0);
 variable VAR_in1 : unsigned(15 downto 0);
 variable VAR_in2 : unsigned(15 downto 0);
 variable VAR_in3 : unsigned(15 downto 0);
 variable VAR_in4 : unsigned(15 downto 0);
 variable VAR_in5 : unsigned(15 downto 0);
 variable VAR_in6 : unsigned(15 downto 0);
 variable VAR_in7 : unsigned(15 downto 0);
 variable VAR_in8 : unsigned(15 downto 0);
 variable VAR_in9 : unsigned(15 downto 0);
 variable VAR_in10 : unsigned(15 downto 0);
 variable VAR_in11 : unsigned(15 downto 0);
 variable VAR_in12 : unsigned(15 downto 0);
 variable VAR_in13 : unsigned(15 downto 0);
 variable VAR_in14 : unsigned(15 downto 0);
 variable VAR_in15 : unsigned(15 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint4_1_1_bit_math_h_l108_c10_4ac4_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint4_2_2_bit_math_h_l158_c10_096f_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_iftrue : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_iffalse : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_iftrue : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_iffalse : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint4_3_3_bit_math_h_l186_c10_0cc5_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iftrue : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iffalse : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_iffalse := VAR_in10;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_iftrue := VAR_in11;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iffalse := VAR_in12;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_iftrue := VAR_in15;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_iffalse := VAR_in2;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_iftrue := VAR_in3;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_iffalse := VAR_in4;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_iftrue := VAR_in5;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_iffalse := VAR_in6;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_iftrue := VAR_in7;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_iffalse := VAR_in8;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_iftrue := VAR_in9;
     -- uint4_0_0[bit_math_h_l14_c10_3c6e] LATENCY=0
     VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output := uint4_0_0(
     VAR_sel);

     -- uint4_3_3[bit_math_h_l186_c10_0cc5] LATENCY=0
     VAR_uint4_3_3_bit_math_h_l186_c10_0cc5_return_output := uint4_3_3(
     VAR_sel);

     -- uint4_2_2[bit_math_h_l158_c10_096f] LATENCY=0
     VAR_uint4_2_2_bit_math_h_l158_c10_096f_return_output := uint4_2_2(
     VAR_sel);

     -- uint4_1_1[bit_math_h_l108_c10_4ac4] LATENCY=0
     VAR_uint4_1_1_bit_math_h_l108_c10_4ac4_return_output := uint4_1_1(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_cond := VAR_uint4_0_0_bit_math_h_l14_c10_3c6e_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_cond := VAR_uint4_1_1_bit_math_h_l108_c10_4ac4_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_cond := VAR_uint4_1_1_bit_math_h_l108_c10_4ac4_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_cond := VAR_uint4_1_1_bit_math_h_l108_c10_4ac4_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_cond := VAR_uint4_1_1_bit_math_h_l108_c10_4ac4_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_cond := VAR_uint4_2_2_bit_math_h_l158_c10_096f_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_cond := VAR_uint4_2_2_bit_math_h_l158_c10_096f_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_cond := VAR_uint4_3_3_bit_math_h_l186_c10_0cc5_return_output;
     -- layer0_node5_MUX[bit_math_h_l73_c3_6697] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_6697_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_6697_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_6697_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output := layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_8dfa] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_8dfa_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output := layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_ee77] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_ee77_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_ee77_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_ee77_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output := layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_d7ea] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_d7ea_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output := layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_c417] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_c417_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_c417_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_c417_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output := layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_55a7] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_55a7_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_55a7_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_55a7_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output := layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_0c13] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_0c13_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_0c13_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_0c13_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output := layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_ee64] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_ee64_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_ee64_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_ee64_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output := layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_8dfa_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_ee77_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_55a7_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_0c13_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_ee64_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_6697_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_d7ea_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_c417_return_output;
     -- layer1_node0_MUX[bit_math_h_l112_c3_a151] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l112_c3_a151_cond <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_cond;
     layer1_node0_MUX_bit_math_h_l112_c3_a151_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_iftrue;
     layer1_node0_MUX_bit_math_h_l112_c3_a151_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output := layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output;

     -- layer1_node2_MUX[bit_math_h_l134_c3_5a40] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l134_c3_5a40_cond <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_cond;
     layer1_node2_MUX_bit_math_h_l134_c3_5a40_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_iftrue;
     layer1_node2_MUX_bit_math_h_l134_c3_5a40_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output := layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output;

     -- layer1_node1_MUX[bit_math_h_l123_c3_f7f1] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l123_c3_f7f1_cond <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_cond;
     layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iftrue;
     layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output := layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output;

     -- layer1_node3_MUX[bit_math_h_l145_c3_b458] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l145_c3_b458_cond <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_cond;
     layer1_node3_MUX_bit_math_h_l145_c3_b458_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_iftrue;
     layer1_node3_MUX_bit_math_h_l145_c3_b458_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output := layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_iffalse := VAR_layer1_node0_MUX_bit_math_h_l112_c3_a151_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_iftrue := VAR_layer1_node1_MUX_bit_math_h_l123_c3_f7f1_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_iffalse := VAR_layer1_node2_MUX_bit_math_h_l134_c3_5a40_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_iftrue := VAR_layer1_node3_MUX_bit_math_h_l145_c3_b458_return_output;
     -- layer2_node1_MUX[bit_math_h_l173_c3_c834] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l173_c3_c834_cond <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_cond;
     layer2_node1_MUX_bit_math_h_l173_c3_c834_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_iftrue;
     layer2_node1_MUX_bit_math_h_l173_c3_c834_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output := layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output;

     -- layer2_node0_MUX[bit_math_h_l162_c3_9803] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l162_c3_9803_cond <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_cond;
     layer2_node0_MUX_bit_math_h_l162_c3_9803_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_iftrue;
     layer2_node0_MUX_bit_math_h_l162_c3_9803_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output := layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iffalse := VAR_layer2_node0_MUX_bit_math_h_l162_c3_9803_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iftrue := VAR_layer2_node1_MUX_bit_math_h_l173_c3_c834_return_output;
     -- layer3_node0_MUX[bit_math_h_l190_c3_d7d1] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l190_c3_d7d1_cond <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_cond;
     layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iftrue;
     layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output := layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output;

     -- Submodule level 5
     VAR_return_output := VAR_layer3_node0_MUX_bit_math_h_l190_c3_d7d1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
